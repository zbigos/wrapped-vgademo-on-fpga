magic
tech sky130A
magscale 1 2
timestamp 1647810391
<< obsli1 >>
rect 1104 527 58880 57681
<< obsm1 >>
rect 566 416 59418 57928
<< metal2 >>
rect 542 59200 654 60000
rect 1646 59200 1758 60000
rect 2842 59200 2954 60000
rect 4038 59200 4150 60000
rect 5234 59200 5346 60000
rect 6338 59200 6450 60000
rect 7534 59200 7646 60000
rect 8730 59200 8842 60000
rect 9926 59200 10038 60000
rect 11122 59200 11234 60000
rect 12226 59200 12338 60000
rect 13422 59200 13534 60000
rect 14618 59200 14730 60000
rect 15814 59200 15926 60000
rect 16918 59200 17030 60000
rect 18114 59200 18226 60000
rect 19310 59200 19422 60000
rect 20506 59200 20618 60000
rect 21702 59200 21814 60000
rect 22806 59200 22918 60000
rect 24002 59200 24114 60000
rect 25198 59200 25310 60000
rect 26394 59200 26506 60000
rect 27590 59200 27702 60000
rect 28694 59200 28806 60000
rect 29890 59200 30002 60000
rect 31086 59200 31198 60000
rect 32282 59200 32394 60000
rect 33386 59200 33498 60000
rect 34582 59200 34694 60000
rect 35778 59200 35890 60000
rect 36974 59200 37086 60000
rect 38170 59200 38282 60000
rect 39274 59200 39386 60000
rect 40470 59200 40582 60000
rect 41666 59200 41778 60000
rect 42862 59200 42974 60000
rect 44058 59200 44170 60000
rect 45162 59200 45274 60000
rect 46358 59200 46470 60000
rect 47554 59200 47666 60000
rect 48750 59200 48862 60000
rect 49854 59200 49966 60000
rect 51050 59200 51162 60000
rect 52246 59200 52358 60000
rect 53442 59200 53554 60000
rect 54638 59200 54750 60000
rect 55742 59200 55854 60000
rect 56938 59200 57050 60000
rect 58134 59200 58246 60000
rect 59330 59200 59442 60000
rect 4222 0 4334 800
rect 12778 0 12890 800
rect 21334 0 21446 800
rect 29890 0 30002 800
rect 38446 0 38558 800
rect 47002 0 47114 800
rect 55558 0 55670 800
<< obsm2 >>
rect 710 59144 1590 59537
rect 1814 59144 2786 59537
rect 3010 59144 3982 59537
rect 4206 59144 5178 59537
rect 5402 59144 6282 59537
rect 6506 59144 7478 59537
rect 7702 59144 8674 59537
rect 8898 59144 9870 59537
rect 10094 59144 11066 59537
rect 11290 59144 12170 59537
rect 12394 59144 13366 59537
rect 13590 59144 14562 59537
rect 14786 59144 15758 59537
rect 15982 59144 16862 59537
rect 17086 59144 18058 59537
rect 18282 59144 19254 59537
rect 19478 59144 20450 59537
rect 20674 59144 21646 59537
rect 21870 59144 22750 59537
rect 22974 59144 23946 59537
rect 24170 59144 25142 59537
rect 25366 59144 26338 59537
rect 26562 59144 27534 59537
rect 27758 59144 28638 59537
rect 28862 59144 29834 59537
rect 30058 59144 31030 59537
rect 31254 59144 32226 59537
rect 32450 59144 33330 59537
rect 33554 59144 34526 59537
rect 34750 59144 35722 59537
rect 35946 59144 36918 59537
rect 37142 59144 38114 59537
rect 38338 59144 39218 59537
rect 39442 59144 40414 59537
rect 40638 59144 41610 59537
rect 41834 59144 42806 59537
rect 43030 59144 44002 59537
rect 44226 59144 45106 59537
rect 45330 59144 46302 59537
rect 46526 59144 47498 59537
rect 47722 59144 48694 59537
rect 48918 59144 49798 59537
rect 50022 59144 50994 59537
rect 51218 59144 52190 59537
rect 52414 59144 53386 59537
rect 53610 59144 54582 59537
rect 54806 59144 55686 59537
rect 55910 59144 56882 59537
rect 57106 59144 58078 59537
rect 58302 59144 59274 59537
rect 572 856 59412 59144
rect 572 410 4166 856
rect 4390 410 12722 856
rect 12946 410 21278 856
rect 21502 410 29834 856
rect 30058 410 38390 856
rect 38614 410 46946 856
rect 47170 410 55502 856
rect 55726 410 59412 856
<< metal3 >>
rect 0 59380 800 59620
rect 59200 59380 60000 59620
rect 0 58564 800 58804
rect 59200 58564 60000 58804
rect 0 57748 800 57988
rect 59200 57884 60000 58124
rect 0 56932 800 57172
rect 59200 57068 60000 57308
rect 0 56116 800 56356
rect 59200 56388 60000 56628
rect 0 55300 800 55540
rect 59200 55572 60000 55812
rect 0 54484 800 54724
rect 59200 54756 60000 54996
rect 59200 54076 60000 54316
rect 0 53668 800 53908
rect 0 52988 800 53228
rect 59200 53260 60000 53500
rect 59200 52580 60000 52820
rect 0 52172 800 52412
rect 59200 51764 60000 52004
rect 0 51356 800 51596
rect 59200 51084 60000 51324
rect 0 50540 800 50780
rect 59200 50268 60000 50508
rect 0 49724 800 49964
rect 59200 49452 60000 49692
rect 0 48908 800 49148
rect 59200 48772 60000 49012
rect 0 48092 800 48332
rect 59200 47956 60000 48196
rect 0 47276 800 47516
rect 59200 47276 60000 47516
rect 0 46596 800 46836
rect 59200 46460 60000 46700
rect 0 45780 800 46020
rect 59200 45644 60000 45884
rect 0 44964 800 45204
rect 59200 44964 60000 45204
rect 0 44148 800 44388
rect 59200 44148 60000 44388
rect 0 43332 800 43572
rect 59200 43468 60000 43708
rect 0 42516 800 42756
rect 59200 42652 60000 42892
rect 0 41700 800 41940
rect 59200 41972 60000 42212
rect 0 40884 800 41124
rect 59200 41156 60000 41396
rect 0 40204 800 40444
rect 59200 40340 60000 40580
rect 0 39388 800 39628
rect 59200 39660 60000 39900
rect 0 38572 800 38812
rect 59200 38844 60000 39084
rect 59200 38164 60000 38404
rect 0 37756 800 37996
rect 59200 37348 60000 37588
rect 0 36940 800 37180
rect 59200 36532 60000 36772
rect 0 36124 800 36364
rect 59200 35852 60000 36092
rect 0 35308 800 35548
rect 59200 35036 60000 35276
rect 0 34492 800 34732
rect 59200 34356 60000 34596
rect 0 33676 800 33916
rect 59200 33540 60000 33780
rect 0 32996 800 33236
rect 59200 32860 60000 33100
rect 0 32180 800 32420
rect 59200 32044 60000 32284
rect 0 31364 800 31604
rect 59200 31228 60000 31468
rect 0 30548 800 30788
rect 59200 30548 60000 30788
rect 0 29732 800 29972
rect 59200 29732 60000 29972
rect 0 28916 800 29156
rect 59200 29052 60000 29292
rect 0 28100 800 28340
rect 59200 28236 60000 28476
rect 0 27284 800 27524
rect 59200 27420 60000 27660
rect 0 26604 800 26844
rect 59200 26740 60000 26980
rect 0 25788 800 26028
rect 59200 25924 60000 26164
rect 0 24972 800 25212
rect 59200 25244 60000 25484
rect 0 24156 800 24396
rect 59200 24428 60000 24668
rect 59200 23748 60000 23988
rect 0 23340 800 23580
rect 59200 22932 60000 23172
rect 0 22524 800 22764
rect 59200 22116 60000 22356
rect 0 21708 800 21948
rect 59200 21436 60000 21676
rect 0 20892 800 21132
rect 59200 20620 60000 20860
rect 0 20212 800 20452
rect 59200 19940 60000 20180
rect 0 19396 800 19636
rect 59200 19124 60000 19364
rect 0 18580 800 18820
rect 59200 18308 60000 18548
rect 0 17764 800 18004
rect 59200 17628 60000 17868
rect 0 16948 800 17188
rect 59200 16812 60000 17052
rect 0 16132 800 16372
rect 59200 16132 60000 16372
rect 0 15316 800 15556
rect 59200 15316 60000 15556
rect 0 14500 800 14740
rect 59200 14636 60000 14876
rect 0 13684 800 13924
rect 59200 13820 60000 14060
rect 0 13004 800 13244
rect 59200 13004 60000 13244
rect 0 12188 800 12428
rect 59200 12324 60000 12564
rect 0 11372 800 11612
rect 59200 11508 60000 11748
rect 0 10556 800 10796
rect 59200 10828 60000 11068
rect 0 9740 800 9980
rect 59200 10012 60000 10252
rect 0 8924 800 9164
rect 59200 9196 60000 9436
rect 59200 8516 60000 8756
rect 0 8108 800 8348
rect 59200 7700 60000 7940
rect 0 7292 800 7532
rect 59200 7020 60000 7260
rect 0 6612 800 6852
rect 59200 6204 60000 6444
rect 0 5796 800 6036
rect 59200 5524 60000 5764
rect 0 4980 800 5220
rect 59200 4708 60000 4948
rect 0 4164 800 4404
rect 59200 3892 60000 4132
rect 0 3348 800 3588
rect 59200 3212 60000 3452
rect 0 2532 800 2772
rect 59200 2396 60000 2636
rect 0 1716 800 1956
rect 59200 1716 60000 1956
rect 0 900 800 1140
rect 59200 900 60000 1140
rect 0 220 800 460
rect 59200 220 60000 460
<< obsm3 >>
rect 880 59300 59120 59533
rect 800 58884 59235 59300
rect 880 58484 59120 58884
rect 800 58204 59235 58484
rect 800 58068 59120 58204
rect 880 57804 59120 58068
rect 880 57668 59235 57804
rect 800 57388 59235 57668
rect 800 57252 59120 57388
rect 880 56988 59120 57252
rect 880 56852 59235 56988
rect 800 56708 59235 56852
rect 800 56436 59120 56708
rect 880 56308 59120 56436
rect 880 56036 59235 56308
rect 800 55892 59235 56036
rect 800 55620 59120 55892
rect 880 55492 59120 55620
rect 880 55220 59235 55492
rect 800 55076 59235 55220
rect 800 54804 59120 55076
rect 880 54676 59120 54804
rect 880 54404 59235 54676
rect 800 54396 59235 54404
rect 800 53996 59120 54396
rect 800 53988 59235 53996
rect 880 53588 59235 53988
rect 800 53580 59235 53588
rect 800 53308 59120 53580
rect 880 53180 59120 53308
rect 880 52908 59235 53180
rect 800 52900 59235 52908
rect 800 52500 59120 52900
rect 800 52492 59235 52500
rect 880 52092 59235 52492
rect 800 52084 59235 52092
rect 800 51684 59120 52084
rect 800 51676 59235 51684
rect 880 51404 59235 51676
rect 880 51276 59120 51404
rect 800 51004 59120 51276
rect 800 50860 59235 51004
rect 880 50588 59235 50860
rect 880 50460 59120 50588
rect 800 50188 59120 50460
rect 800 50044 59235 50188
rect 880 49772 59235 50044
rect 880 49644 59120 49772
rect 800 49372 59120 49644
rect 800 49228 59235 49372
rect 880 49092 59235 49228
rect 880 48828 59120 49092
rect 800 48692 59120 48828
rect 800 48412 59235 48692
rect 880 48276 59235 48412
rect 880 48012 59120 48276
rect 800 47876 59120 48012
rect 800 47596 59235 47876
rect 880 47196 59120 47596
rect 800 46916 59235 47196
rect 880 46780 59235 46916
rect 880 46516 59120 46780
rect 800 46380 59120 46516
rect 800 46100 59235 46380
rect 880 45964 59235 46100
rect 880 45700 59120 45964
rect 800 45564 59120 45700
rect 800 45284 59235 45564
rect 880 44884 59120 45284
rect 800 44468 59235 44884
rect 880 44068 59120 44468
rect 800 43788 59235 44068
rect 800 43652 59120 43788
rect 880 43388 59120 43652
rect 880 43252 59235 43388
rect 800 42972 59235 43252
rect 800 42836 59120 42972
rect 880 42572 59120 42836
rect 880 42436 59235 42572
rect 800 42292 59235 42436
rect 800 42020 59120 42292
rect 880 41892 59120 42020
rect 880 41620 59235 41892
rect 800 41476 59235 41620
rect 800 41204 59120 41476
rect 880 41076 59120 41204
rect 880 40804 59235 41076
rect 800 40660 59235 40804
rect 800 40524 59120 40660
rect 880 40260 59120 40524
rect 880 40124 59235 40260
rect 800 39980 59235 40124
rect 800 39708 59120 39980
rect 880 39580 59120 39708
rect 880 39308 59235 39580
rect 800 39164 59235 39308
rect 800 38892 59120 39164
rect 880 38764 59120 38892
rect 880 38492 59235 38764
rect 800 38484 59235 38492
rect 800 38084 59120 38484
rect 800 38076 59235 38084
rect 880 37676 59235 38076
rect 800 37668 59235 37676
rect 800 37268 59120 37668
rect 800 37260 59235 37268
rect 880 36860 59235 37260
rect 800 36852 59235 36860
rect 800 36452 59120 36852
rect 800 36444 59235 36452
rect 880 36172 59235 36444
rect 880 36044 59120 36172
rect 800 35772 59120 36044
rect 800 35628 59235 35772
rect 880 35356 59235 35628
rect 880 35228 59120 35356
rect 800 34956 59120 35228
rect 800 34812 59235 34956
rect 880 34676 59235 34812
rect 880 34412 59120 34676
rect 800 34276 59120 34412
rect 800 33996 59235 34276
rect 880 33860 59235 33996
rect 880 33596 59120 33860
rect 800 33460 59120 33596
rect 800 33316 59235 33460
rect 880 33180 59235 33316
rect 880 32916 59120 33180
rect 800 32780 59120 32916
rect 800 32500 59235 32780
rect 880 32364 59235 32500
rect 880 32100 59120 32364
rect 800 31964 59120 32100
rect 800 31684 59235 31964
rect 880 31548 59235 31684
rect 880 31284 59120 31548
rect 800 31148 59120 31284
rect 800 30868 59235 31148
rect 880 30468 59120 30868
rect 800 30052 59235 30468
rect 880 29652 59120 30052
rect 800 29372 59235 29652
rect 800 29236 59120 29372
rect 880 28972 59120 29236
rect 880 28836 59235 28972
rect 800 28556 59235 28836
rect 800 28420 59120 28556
rect 880 28156 59120 28420
rect 880 28020 59235 28156
rect 800 27740 59235 28020
rect 800 27604 59120 27740
rect 880 27340 59120 27604
rect 880 27204 59235 27340
rect 800 27060 59235 27204
rect 800 26924 59120 27060
rect 880 26660 59120 26924
rect 880 26524 59235 26660
rect 800 26244 59235 26524
rect 800 26108 59120 26244
rect 880 25844 59120 26108
rect 880 25708 59235 25844
rect 800 25564 59235 25708
rect 800 25292 59120 25564
rect 880 25164 59120 25292
rect 880 24892 59235 25164
rect 800 24748 59235 24892
rect 800 24476 59120 24748
rect 880 24348 59120 24476
rect 880 24076 59235 24348
rect 800 24068 59235 24076
rect 800 23668 59120 24068
rect 800 23660 59235 23668
rect 880 23260 59235 23660
rect 800 23252 59235 23260
rect 800 22852 59120 23252
rect 800 22844 59235 22852
rect 880 22444 59235 22844
rect 800 22436 59235 22444
rect 800 22036 59120 22436
rect 800 22028 59235 22036
rect 880 21756 59235 22028
rect 880 21628 59120 21756
rect 800 21356 59120 21628
rect 800 21212 59235 21356
rect 880 20940 59235 21212
rect 880 20812 59120 20940
rect 800 20540 59120 20812
rect 800 20532 59235 20540
rect 880 20260 59235 20532
rect 880 20132 59120 20260
rect 800 19860 59120 20132
rect 800 19716 59235 19860
rect 880 19444 59235 19716
rect 880 19316 59120 19444
rect 800 19044 59120 19316
rect 800 18900 59235 19044
rect 880 18628 59235 18900
rect 880 18500 59120 18628
rect 800 18228 59120 18500
rect 800 18084 59235 18228
rect 880 17948 59235 18084
rect 880 17684 59120 17948
rect 800 17548 59120 17684
rect 800 17268 59235 17548
rect 880 17132 59235 17268
rect 880 16868 59120 17132
rect 800 16732 59120 16868
rect 800 16452 59235 16732
rect 880 16052 59120 16452
rect 800 15636 59235 16052
rect 880 15236 59120 15636
rect 800 14956 59235 15236
rect 800 14820 59120 14956
rect 880 14556 59120 14820
rect 880 14420 59235 14556
rect 800 14140 59235 14420
rect 800 14004 59120 14140
rect 880 13740 59120 14004
rect 880 13604 59235 13740
rect 800 13324 59235 13604
rect 880 12924 59120 13324
rect 800 12644 59235 12924
rect 800 12508 59120 12644
rect 880 12244 59120 12508
rect 880 12108 59235 12244
rect 800 11828 59235 12108
rect 800 11692 59120 11828
rect 880 11428 59120 11692
rect 880 11292 59235 11428
rect 800 11148 59235 11292
rect 800 10876 59120 11148
rect 880 10748 59120 10876
rect 880 10476 59235 10748
rect 800 10332 59235 10476
rect 800 10060 59120 10332
rect 880 9932 59120 10060
rect 880 9660 59235 9932
rect 800 9516 59235 9660
rect 800 9244 59120 9516
rect 880 9116 59120 9244
rect 880 8844 59235 9116
rect 800 8836 59235 8844
rect 800 8436 59120 8836
rect 800 8428 59235 8436
rect 880 8028 59235 8428
rect 800 8020 59235 8028
rect 800 7620 59120 8020
rect 800 7612 59235 7620
rect 880 7340 59235 7612
rect 880 7212 59120 7340
rect 800 6940 59120 7212
rect 800 6932 59235 6940
rect 880 6532 59235 6932
rect 800 6524 59235 6532
rect 800 6124 59120 6524
rect 800 6116 59235 6124
rect 880 5844 59235 6116
rect 880 5716 59120 5844
rect 800 5444 59120 5716
rect 800 5300 59235 5444
rect 880 5028 59235 5300
rect 880 4900 59120 5028
rect 800 4628 59120 4900
rect 800 4484 59235 4628
rect 880 4212 59235 4484
rect 880 4084 59120 4212
rect 800 3812 59120 4084
rect 800 3668 59235 3812
rect 880 3532 59235 3668
rect 880 3268 59120 3532
rect 800 3132 59120 3268
rect 800 2852 59235 3132
rect 880 2716 59235 2852
rect 880 2452 59120 2716
rect 800 2316 59120 2452
rect 800 2036 59235 2316
rect 880 1636 59120 2036
rect 800 1220 59235 1636
rect 880 820 59120 1220
rect 800 540 59235 820
rect 880 511 59120 540
<< metal4 >>
rect 4208 496 4528 57712
rect 19568 496 19888 57712
rect 34928 496 35248 57712
rect 50288 496 50608 57712
<< obsm4 >>
rect 19195 3435 19488 54365
rect 19968 3435 34848 54365
rect 35328 3435 50208 54365
rect 50688 3435 57717 54365
<< labels >>
rlabel metal2 s 542 59200 654 60000 6 active
port 1 nsew signal input
rlabel metal2 s 2842 59200 2954 60000 6 io_in[0]
port 2 nsew signal input
rlabel metal2 s 14618 59200 14730 60000 6 io_in[10]
port 3 nsew signal input
rlabel metal2 s 15814 59200 15926 60000 6 io_in[11]
port 4 nsew signal input
rlabel metal2 s 16918 59200 17030 60000 6 io_in[12]
port 5 nsew signal input
rlabel metal2 s 18114 59200 18226 60000 6 io_in[13]
port 6 nsew signal input
rlabel metal2 s 19310 59200 19422 60000 6 io_in[14]
port 7 nsew signal input
rlabel metal2 s 20506 59200 20618 60000 6 io_in[15]
port 8 nsew signal input
rlabel metal2 s 21702 59200 21814 60000 6 io_in[16]
port 9 nsew signal input
rlabel metal2 s 22806 59200 22918 60000 6 io_in[17]
port 10 nsew signal input
rlabel metal2 s 24002 59200 24114 60000 6 io_in[18]
port 11 nsew signal input
rlabel metal2 s 25198 59200 25310 60000 6 io_in[19]
port 12 nsew signal input
rlabel metal2 s 4038 59200 4150 60000 6 io_in[1]
port 13 nsew signal input
rlabel metal2 s 26394 59200 26506 60000 6 io_in[20]
port 14 nsew signal input
rlabel metal2 s 27590 59200 27702 60000 6 io_in[21]
port 15 nsew signal input
rlabel metal2 s 28694 59200 28806 60000 6 io_in[22]
port 16 nsew signal input
rlabel metal2 s 29890 59200 30002 60000 6 io_in[23]
port 17 nsew signal input
rlabel metal2 s 31086 59200 31198 60000 6 io_in[24]
port 18 nsew signal input
rlabel metal2 s 32282 59200 32394 60000 6 io_in[25]
port 19 nsew signal input
rlabel metal2 s 33386 59200 33498 60000 6 io_in[26]
port 20 nsew signal input
rlabel metal2 s 34582 59200 34694 60000 6 io_in[27]
port 21 nsew signal input
rlabel metal2 s 35778 59200 35890 60000 6 io_in[28]
port 22 nsew signal input
rlabel metal2 s 36974 59200 37086 60000 6 io_in[29]
port 23 nsew signal input
rlabel metal2 s 5234 59200 5346 60000 6 io_in[2]
port 24 nsew signal input
rlabel metal2 s 38170 59200 38282 60000 6 io_in[30]
port 25 nsew signal input
rlabel metal2 s 39274 59200 39386 60000 6 io_in[31]
port 26 nsew signal input
rlabel metal2 s 40470 59200 40582 60000 6 io_in[32]
port 27 nsew signal input
rlabel metal2 s 41666 59200 41778 60000 6 io_in[33]
port 28 nsew signal input
rlabel metal2 s 42862 59200 42974 60000 6 io_in[34]
port 29 nsew signal input
rlabel metal2 s 44058 59200 44170 60000 6 io_in[35]
port 30 nsew signal input
rlabel metal2 s 45162 59200 45274 60000 6 io_in[36]
port 31 nsew signal input
rlabel metal2 s 46358 59200 46470 60000 6 io_in[37]
port 32 nsew signal input
rlabel metal2 s 6338 59200 6450 60000 6 io_in[3]
port 33 nsew signal input
rlabel metal2 s 7534 59200 7646 60000 6 io_in[4]
port 34 nsew signal input
rlabel metal2 s 8730 59200 8842 60000 6 io_in[5]
port 35 nsew signal input
rlabel metal2 s 9926 59200 10038 60000 6 io_in[6]
port 36 nsew signal input
rlabel metal2 s 11122 59200 11234 60000 6 io_in[7]
port 37 nsew signal input
rlabel metal2 s 12226 59200 12338 60000 6 io_in[8]
port 38 nsew signal input
rlabel metal2 s 13422 59200 13534 60000 6 io_in[9]
port 39 nsew signal input
rlabel metal3 s 59200 24428 60000 24668 6 io_oeb[0]
port 40 nsew signal output
rlabel metal3 s 59200 32044 60000 32284 6 io_oeb[10]
port 41 nsew signal output
rlabel metal3 s 59200 32860 60000 33100 6 io_oeb[11]
port 42 nsew signal output
rlabel metal3 s 59200 33540 60000 33780 6 io_oeb[12]
port 43 nsew signal output
rlabel metal3 s 59200 34356 60000 34596 6 io_oeb[13]
port 44 nsew signal output
rlabel metal3 s 59200 35036 60000 35276 6 io_oeb[14]
port 45 nsew signal output
rlabel metal3 s 59200 35852 60000 36092 6 io_oeb[15]
port 46 nsew signal output
rlabel metal3 s 59200 36532 60000 36772 6 io_oeb[16]
port 47 nsew signal output
rlabel metal3 s 59200 37348 60000 37588 6 io_oeb[17]
port 48 nsew signal output
rlabel metal3 s 59200 38164 60000 38404 6 io_oeb[18]
port 49 nsew signal output
rlabel metal3 s 59200 38844 60000 39084 6 io_oeb[19]
port 50 nsew signal output
rlabel metal3 s 59200 25244 60000 25484 6 io_oeb[1]
port 51 nsew signal output
rlabel metal3 s 59200 39660 60000 39900 6 io_oeb[20]
port 52 nsew signal output
rlabel metal3 s 59200 40340 60000 40580 6 io_oeb[21]
port 53 nsew signal output
rlabel metal3 s 59200 41156 60000 41396 6 io_oeb[22]
port 54 nsew signal output
rlabel metal3 s 59200 41972 60000 42212 6 io_oeb[23]
port 55 nsew signal output
rlabel metal3 s 59200 42652 60000 42892 6 io_oeb[24]
port 56 nsew signal output
rlabel metal3 s 59200 43468 60000 43708 6 io_oeb[25]
port 57 nsew signal output
rlabel metal3 s 59200 44148 60000 44388 6 io_oeb[26]
port 58 nsew signal output
rlabel metal3 s 59200 44964 60000 45204 6 io_oeb[27]
port 59 nsew signal output
rlabel metal3 s 59200 45644 60000 45884 6 io_oeb[28]
port 60 nsew signal output
rlabel metal3 s 59200 46460 60000 46700 6 io_oeb[29]
port 61 nsew signal output
rlabel metal3 s 59200 25924 60000 26164 6 io_oeb[2]
port 62 nsew signal output
rlabel metal3 s 59200 47276 60000 47516 6 io_oeb[30]
port 63 nsew signal output
rlabel metal3 s 59200 47956 60000 48196 6 io_oeb[31]
port 64 nsew signal output
rlabel metal3 s 59200 48772 60000 49012 6 io_oeb[32]
port 65 nsew signal output
rlabel metal3 s 59200 49452 60000 49692 6 io_oeb[33]
port 66 nsew signal output
rlabel metal3 s 59200 50268 60000 50508 6 io_oeb[34]
port 67 nsew signal output
rlabel metal3 s 59200 51084 60000 51324 6 io_oeb[35]
port 68 nsew signal output
rlabel metal3 s 59200 51764 60000 52004 6 io_oeb[36]
port 69 nsew signal output
rlabel metal3 s 59200 52580 60000 52820 6 io_oeb[37]
port 70 nsew signal output
rlabel metal3 s 59200 26740 60000 26980 6 io_oeb[3]
port 71 nsew signal output
rlabel metal3 s 59200 27420 60000 27660 6 io_oeb[4]
port 72 nsew signal output
rlabel metal3 s 59200 28236 60000 28476 6 io_oeb[5]
port 73 nsew signal output
rlabel metal3 s 59200 29052 60000 29292 6 io_oeb[6]
port 74 nsew signal output
rlabel metal3 s 59200 29732 60000 29972 6 io_oeb[7]
port 75 nsew signal output
rlabel metal3 s 59200 30548 60000 30788 6 io_oeb[8]
port 76 nsew signal output
rlabel metal3 s 59200 31228 60000 31468 6 io_oeb[9]
port 77 nsew signal output
rlabel metal3 s 59200 53260 60000 53500 6 io_out[0]
port 78 nsew signal output
rlabel metal3 s 0 53668 800 53908 6 io_out[10]
port 79 nsew signal output
rlabel metal3 s 59200 55572 60000 55812 6 io_out[11]
port 80 nsew signal output
rlabel metal3 s 59200 56388 60000 56628 6 io_out[12]
port 81 nsew signal output
rlabel metal3 s 59200 57068 60000 57308 6 io_out[13]
port 82 nsew signal output
rlabel metal2 s 12778 0 12890 800 6 io_out[14]
port 83 nsew signal output
rlabel metal2 s 51050 59200 51162 60000 6 io_out[15]
port 84 nsew signal output
rlabel metal3 s 0 54484 800 54724 6 io_out[16]
port 85 nsew signal output
rlabel metal3 s 59200 57884 60000 58124 6 io_out[17]
port 86 nsew signal output
rlabel metal2 s 52246 59200 52358 60000 6 io_out[18]
port 87 nsew signal output
rlabel metal2 s 53442 59200 53554 60000 6 io_out[19]
port 88 nsew signal output
rlabel metal3 s 59200 54076 60000 54316 6 io_out[1]
port 89 nsew signal output
rlabel metal2 s 54638 59200 54750 60000 6 io_out[20]
port 90 nsew signal output
rlabel metal2 s 21334 0 21446 800 6 io_out[21]
port 91 nsew signal output
rlabel metal3 s 0 55300 800 55540 6 io_out[22]
port 92 nsew signal output
rlabel metal2 s 29890 0 30002 800 6 io_out[23]
port 93 nsew signal output
rlabel metal2 s 55742 59200 55854 60000 6 io_out[24]
port 94 nsew signal output
rlabel metal3 s 59200 58564 60000 58804 6 io_out[25]
port 95 nsew signal output
rlabel metal3 s 0 56116 800 56356 6 io_out[26]
port 96 nsew signal output
rlabel metal2 s 38446 0 38558 800 6 io_out[27]
port 97 nsew signal output
rlabel metal2 s 47002 0 47114 800 6 io_out[28]
port 98 nsew signal output
rlabel metal3 s 59200 59380 60000 59620 6 io_out[29]
port 99 nsew signal output
rlabel metal3 s 0 51356 800 51596 6 io_out[2]
port 100 nsew signal output
rlabel metal2 s 56938 59200 57050 60000 6 io_out[30]
port 101 nsew signal output
rlabel metal2 s 58134 59200 58246 60000 6 io_out[31]
port 102 nsew signal output
rlabel metal3 s 0 56932 800 57172 6 io_out[32]
port 103 nsew signal output
rlabel metal3 s 0 57748 800 57988 6 io_out[33]
port 104 nsew signal output
rlabel metal3 s 0 58564 800 58804 6 io_out[34]
port 105 nsew signal output
rlabel metal2 s 59330 59200 59442 60000 6 io_out[35]
port 106 nsew signal output
rlabel metal3 s 0 59380 800 59620 6 io_out[36]
port 107 nsew signal output
rlabel metal2 s 55558 0 55670 800 6 io_out[37]
port 108 nsew signal output
rlabel metal3 s 0 52172 800 52412 6 io_out[3]
port 109 nsew signal output
rlabel metal2 s 47554 59200 47666 60000 6 io_out[4]
port 110 nsew signal output
rlabel metal3 s 0 52988 800 53228 6 io_out[5]
port 111 nsew signal output
rlabel metal2 s 48750 59200 48862 60000 6 io_out[6]
port 112 nsew signal output
rlabel metal2 s 49854 59200 49966 60000 6 io_out[7]
port 113 nsew signal output
rlabel metal2 s 4222 0 4334 800 6 io_out[8]
port 114 nsew signal output
rlabel metal3 s 59200 54756 60000 54996 6 io_out[9]
port 115 nsew signal output
rlabel metal3 s 0 220 800 460 6 la1_data_in[0]
port 116 nsew signal input
rlabel metal3 s 0 8108 800 8348 6 la1_data_in[10]
port 117 nsew signal input
rlabel metal3 s 0 8924 800 9164 6 la1_data_in[11]
port 118 nsew signal input
rlabel metal3 s 0 9740 800 9980 6 la1_data_in[12]
port 119 nsew signal input
rlabel metal3 s 0 10556 800 10796 6 la1_data_in[13]
port 120 nsew signal input
rlabel metal3 s 0 11372 800 11612 6 la1_data_in[14]
port 121 nsew signal input
rlabel metal3 s 0 12188 800 12428 6 la1_data_in[15]
port 122 nsew signal input
rlabel metal3 s 0 13004 800 13244 6 la1_data_in[16]
port 123 nsew signal input
rlabel metal3 s 0 13684 800 13924 6 la1_data_in[17]
port 124 nsew signal input
rlabel metal3 s 0 14500 800 14740 6 la1_data_in[18]
port 125 nsew signal input
rlabel metal3 s 0 15316 800 15556 6 la1_data_in[19]
port 126 nsew signal input
rlabel metal3 s 0 900 800 1140 6 la1_data_in[1]
port 127 nsew signal input
rlabel metal3 s 0 16132 800 16372 6 la1_data_in[20]
port 128 nsew signal input
rlabel metal3 s 0 16948 800 17188 6 la1_data_in[21]
port 129 nsew signal input
rlabel metal3 s 0 17764 800 18004 6 la1_data_in[22]
port 130 nsew signal input
rlabel metal3 s 0 18580 800 18820 6 la1_data_in[23]
port 131 nsew signal input
rlabel metal3 s 0 19396 800 19636 6 la1_data_in[24]
port 132 nsew signal input
rlabel metal3 s 0 20212 800 20452 6 la1_data_in[25]
port 133 nsew signal input
rlabel metal3 s 0 20892 800 21132 6 la1_data_in[26]
port 134 nsew signal input
rlabel metal3 s 0 21708 800 21948 6 la1_data_in[27]
port 135 nsew signal input
rlabel metal3 s 0 22524 800 22764 6 la1_data_in[28]
port 136 nsew signal input
rlabel metal3 s 0 23340 800 23580 6 la1_data_in[29]
port 137 nsew signal input
rlabel metal3 s 0 1716 800 1956 6 la1_data_in[2]
port 138 nsew signal input
rlabel metal3 s 0 24156 800 24396 6 la1_data_in[30]
port 139 nsew signal input
rlabel metal3 s 0 24972 800 25212 6 la1_data_in[31]
port 140 nsew signal input
rlabel metal3 s 0 2532 800 2772 6 la1_data_in[3]
port 141 nsew signal input
rlabel metal3 s 0 3348 800 3588 6 la1_data_in[4]
port 142 nsew signal input
rlabel metal3 s 0 4164 800 4404 6 la1_data_in[5]
port 143 nsew signal input
rlabel metal3 s 0 4980 800 5220 6 la1_data_in[6]
port 144 nsew signal input
rlabel metal3 s 0 5796 800 6036 6 la1_data_in[7]
port 145 nsew signal input
rlabel metal3 s 0 6612 800 6852 6 la1_data_in[8]
port 146 nsew signal input
rlabel metal3 s 0 7292 800 7532 6 la1_data_in[9]
port 147 nsew signal input
rlabel metal3 s 0 25788 800 26028 6 la1_data_out[0]
port 148 nsew signal output
rlabel metal3 s 0 33676 800 33916 6 la1_data_out[10]
port 149 nsew signal output
rlabel metal3 s 0 34492 800 34732 6 la1_data_out[11]
port 150 nsew signal output
rlabel metal3 s 0 35308 800 35548 6 la1_data_out[12]
port 151 nsew signal output
rlabel metal3 s 0 36124 800 36364 6 la1_data_out[13]
port 152 nsew signal output
rlabel metal3 s 0 36940 800 37180 6 la1_data_out[14]
port 153 nsew signal output
rlabel metal3 s 0 37756 800 37996 6 la1_data_out[15]
port 154 nsew signal output
rlabel metal3 s 0 38572 800 38812 6 la1_data_out[16]
port 155 nsew signal output
rlabel metal3 s 0 39388 800 39628 6 la1_data_out[17]
port 156 nsew signal output
rlabel metal3 s 0 40204 800 40444 6 la1_data_out[18]
port 157 nsew signal output
rlabel metal3 s 0 40884 800 41124 6 la1_data_out[19]
port 158 nsew signal output
rlabel metal3 s 0 26604 800 26844 6 la1_data_out[1]
port 159 nsew signal output
rlabel metal3 s 0 41700 800 41940 6 la1_data_out[20]
port 160 nsew signal output
rlabel metal3 s 0 42516 800 42756 6 la1_data_out[21]
port 161 nsew signal output
rlabel metal3 s 0 43332 800 43572 6 la1_data_out[22]
port 162 nsew signal output
rlabel metal3 s 0 44148 800 44388 6 la1_data_out[23]
port 163 nsew signal output
rlabel metal3 s 0 44964 800 45204 6 la1_data_out[24]
port 164 nsew signal output
rlabel metal3 s 0 45780 800 46020 6 la1_data_out[25]
port 165 nsew signal output
rlabel metal3 s 0 46596 800 46836 6 la1_data_out[26]
port 166 nsew signal output
rlabel metal3 s 0 47276 800 47516 6 la1_data_out[27]
port 167 nsew signal output
rlabel metal3 s 0 48092 800 48332 6 la1_data_out[28]
port 168 nsew signal output
rlabel metal3 s 0 48908 800 49148 6 la1_data_out[29]
port 169 nsew signal output
rlabel metal3 s 0 27284 800 27524 6 la1_data_out[2]
port 170 nsew signal output
rlabel metal3 s 0 49724 800 49964 6 la1_data_out[30]
port 171 nsew signal output
rlabel metal3 s 0 50540 800 50780 6 la1_data_out[31]
port 172 nsew signal output
rlabel metal3 s 0 28100 800 28340 6 la1_data_out[3]
port 173 nsew signal output
rlabel metal3 s 0 28916 800 29156 6 la1_data_out[4]
port 174 nsew signal output
rlabel metal3 s 0 29732 800 29972 6 la1_data_out[5]
port 175 nsew signal output
rlabel metal3 s 0 30548 800 30788 6 la1_data_out[6]
port 176 nsew signal output
rlabel metal3 s 0 31364 800 31604 6 la1_data_out[7]
port 177 nsew signal output
rlabel metal3 s 0 32180 800 32420 6 la1_data_out[8]
port 178 nsew signal output
rlabel metal3 s 0 32996 800 33236 6 la1_data_out[9]
port 179 nsew signal output
rlabel metal3 s 59200 220 60000 460 6 la1_oenb[0]
port 180 nsew signal input
rlabel metal3 s 59200 7700 60000 7940 6 la1_oenb[10]
port 181 nsew signal input
rlabel metal3 s 59200 8516 60000 8756 6 la1_oenb[11]
port 182 nsew signal input
rlabel metal3 s 59200 9196 60000 9436 6 la1_oenb[12]
port 183 nsew signal input
rlabel metal3 s 59200 10012 60000 10252 6 la1_oenb[13]
port 184 nsew signal input
rlabel metal3 s 59200 10828 60000 11068 6 la1_oenb[14]
port 185 nsew signal input
rlabel metal3 s 59200 11508 60000 11748 6 la1_oenb[15]
port 186 nsew signal input
rlabel metal3 s 59200 12324 60000 12564 6 la1_oenb[16]
port 187 nsew signal input
rlabel metal3 s 59200 13004 60000 13244 6 la1_oenb[17]
port 188 nsew signal input
rlabel metal3 s 59200 13820 60000 14060 6 la1_oenb[18]
port 189 nsew signal input
rlabel metal3 s 59200 14636 60000 14876 6 la1_oenb[19]
port 190 nsew signal input
rlabel metal3 s 59200 900 60000 1140 6 la1_oenb[1]
port 191 nsew signal input
rlabel metal3 s 59200 15316 60000 15556 6 la1_oenb[20]
port 192 nsew signal input
rlabel metal3 s 59200 16132 60000 16372 6 la1_oenb[21]
port 193 nsew signal input
rlabel metal3 s 59200 16812 60000 17052 6 la1_oenb[22]
port 194 nsew signal input
rlabel metal3 s 59200 17628 60000 17868 6 la1_oenb[23]
port 195 nsew signal input
rlabel metal3 s 59200 18308 60000 18548 6 la1_oenb[24]
port 196 nsew signal input
rlabel metal3 s 59200 19124 60000 19364 6 la1_oenb[25]
port 197 nsew signal input
rlabel metal3 s 59200 19940 60000 20180 6 la1_oenb[26]
port 198 nsew signal input
rlabel metal3 s 59200 20620 60000 20860 6 la1_oenb[27]
port 199 nsew signal input
rlabel metal3 s 59200 21436 60000 21676 6 la1_oenb[28]
port 200 nsew signal input
rlabel metal3 s 59200 22116 60000 22356 6 la1_oenb[29]
port 201 nsew signal input
rlabel metal3 s 59200 1716 60000 1956 6 la1_oenb[2]
port 202 nsew signal input
rlabel metal3 s 59200 22932 60000 23172 6 la1_oenb[30]
port 203 nsew signal input
rlabel metal3 s 59200 23748 60000 23988 6 la1_oenb[31]
port 204 nsew signal input
rlabel metal3 s 59200 2396 60000 2636 6 la1_oenb[3]
port 205 nsew signal input
rlabel metal3 s 59200 3212 60000 3452 6 la1_oenb[4]
port 206 nsew signal input
rlabel metal3 s 59200 3892 60000 4132 6 la1_oenb[5]
port 207 nsew signal input
rlabel metal3 s 59200 4708 60000 4948 6 la1_oenb[6]
port 208 nsew signal input
rlabel metal3 s 59200 5524 60000 5764 6 la1_oenb[7]
port 209 nsew signal input
rlabel metal3 s 59200 6204 60000 6444 6 la1_oenb[8]
port 210 nsew signal input
rlabel metal3 s 59200 7020 60000 7260 6 la1_oenb[9]
port 211 nsew signal input
rlabel metal4 s 4208 496 4528 57712 6 vccd1
port 212 nsew power input
rlabel metal4 s 34928 496 35248 57712 6 vccd1
port 212 nsew power input
rlabel metal4 s 19568 496 19888 57712 6 vssd1
port 213 nsew ground input
rlabel metal4 s 50288 496 50608 57712 6 vssd1
port 213 nsew ground input
rlabel metal2 s 1646 59200 1758 60000 6 wb_clk_i
port 214 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 60000 60000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 12668874
string GDS_FILE /openlane/designs/wrapped-vgademo-on-fpga/runs/RUN_2022.03.20_21.01.03/results/finishing/wrapped_vgademo_on_fpga.magic.gds
string GDS_START 1072870
<< end >>

