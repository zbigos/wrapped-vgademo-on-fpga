magic
tech sky130A
magscale 1 2
timestamp 1647762466
<< obsli1 >>
rect 1104 527 58880 57681
<< obsm1 >>
rect 566 280 59418 57792
<< metal2 >>
rect 542 59200 654 60000
rect 1646 59200 1758 60000
rect 2750 59200 2862 60000
rect 3854 59200 3966 60000
rect 5050 59200 5162 60000
rect 6154 59200 6266 60000
rect 7258 59200 7370 60000
rect 8454 59200 8566 60000
rect 9558 59200 9670 60000
rect 10662 59200 10774 60000
rect 11858 59200 11970 60000
rect 12962 59200 13074 60000
rect 14066 59200 14178 60000
rect 15170 59200 15282 60000
rect 16366 59200 16478 60000
rect 17470 59200 17582 60000
rect 18574 59200 18686 60000
rect 19770 59200 19882 60000
rect 20874 59200 20986 60000
rect 21978 59200 22090 60000
rect 23174 59200 23286 60000
rect 24278 59200 24390 60000
rect 25382 59200 25494 60000
rect 26486 59200 26598 60000
rect 27682 59200 27794 60000
rect 28786 59200 28898 60000
rect 29890 59200 30002 60000
rect 31086 59200 31198 60000
rect 32190 59200 32302 60000
rect 33294 59200 33406 60000
rect 34490 59200 34602 60000
rect 35594 59200 35706 60000
rect 36698 59200 36810 60000
rect 37802 59200 37914 60000
rect 38998 59200 39110 60000
rect 40102 59200 40214 60000
rect 41206 59200 41318 60000
rect 42402 59200 42514 60000
rect 43506 59200 43618 60000
rect 44610 59200 44722 60000
rect 45806 59200 45918 60000
rect 46910 59200 47022 60000
rect 48014 59200 48126 60000
rect 49118 59200 49230 60000
rect 50314 59200 50426 60000
rect 51418 59200 51530 60000
rect 52522 59200 52634 60000
rect 53718 59200 53830 60000
rect 54822 59200 54934 60000
rect 55926 59200 56038 60000
rect 57122 59200 57234 60000
rect 58226 59200 58338 60000
rect 59330 59200 59442 60000
rect 3670 0 3782 800
rect 11122 0 11234 800
rect 18666 0 18778 800
rect 26118 0 26230 800
rect 33662 0 33774 800
rect 41114 0 41226 800
rect 48658 0 48770 800
rect 56110 0 56222 800
<< obsm2 >>
rect 710 59144 1590 59537
rect 1814 59144 2694 59537
rect 2918 59144 3798 59537
rect 4022 59144 4994 59537
rect 5218 59144 6098 59537
rect 6322 59144 7202 59537
rect 7426 59144 8398 59537
rect 8622 59144 9502 59537
rect 9726 59144 10606 59537
rect 10830 59144 11802 59537
rect 12026 59144 12906 59537
rect 13130 59144 14010 59537
rect 14234 59144 15114 59537
rect 15338 59144 16310 59537
rect 16534 59144 17414 59537
rect 17638 59144 18518 59537
rect 18742 59144 19714 59537
rect 19938 59144 20818 59537
rect 21042 59144 21922 59537
rect 22146 59144 23118 59537
rect 23342 59144 24222 59537
rect 24446 59144 25326 59537
rect 25550 59144 26430 59537
rect 26654 59144 27626 59537
rect 27850 59144 28730 59537
rect 28954 59144 29834 59537
rect 30058 59144 31030 59537
rect 31254 59144 32134 59537
rect 32358 59144 33238 59537
rect 33462 59144 34434 59537
rect 34658 59144 35538 59537
rect 35762 59144 36642 59537
rect 36866 59144 37746 59537
rect 37970 59144 38942 59537
rect 39166 59144 40046 59537
rect 40270 59144 41150 59537
rect 41374 59144 42346 59537
rect 42570 59144 43450 59537
rect 43674 59144 44554 59537
rect 44778 59144 45750 59537
rect 45974 59144 46854 59537
rect 47078 59144 47958 59537
rect 48182 59144 49062 59537
rect 49286 59144 50258 59537
rect 50482 59144 51362 59537
rect 51586 59144 52466 59537
rect 52690 59144 53662 59537
rect 53886 59144 54766 59537
rect 54990 59144 55870 59537
rect 56094 59144 57066 59537
rect 57290 59144 58170 59537
rect 58394 59144 59274 59537
rect 572 856 59412 59144
rect 572 274 3614 856
rect 3838 274 11066 856
rect 11290 274 18610 856
rect 18834 274 26062 856
rect 26286 274 33606 856
rect 33830 274 41058 856
rect 41282 274 48602 856
rect 48826 274 56054 856
rect 56278 274 59412 856
<< metal3 >>
rect 0 59380 800 59620
rect 59200 59380 60000 59620
rect 0 58564 800 58804
rect 59200 58564 60000 58804
rect 0 57748 800 57988
rect 59200 57884 60000 58124
rect 0 56932 800 57172
rect 59200 57068 60000 57308
rect 0 56116 800 56356
rect 59200 56388 60000 56628
rect 0 55300 800 55540
rect 59200 55572 60000 55812
rect 0 54484 800 54724
rect 59200 54756 60000 54996
rect 59200 54076 60000 54316
rect 0 53668 800 53908
rect 59200 53260 60000 53500
rect 0 52716 800 52956
rect 59200 52580 60000 52820
rect 0 51900 800 52140
rect 59200 51764 60000 52004
rect 0 51084 800 51324
rect 59200 51084 60000 51324
rect 0 50268 800 50508
rect 59200 50268 60000 50508
rect 0 49452 800 49692
rect 59200 49452 60000 49692
rect 0 48636 800 48876
rect 59200 48772 60000 49012
rect 0 47820 800 48060
rect 59200 47956 60000 48196
rect 0 47004 800 47244
rect 59200 47276 60000 47516
rect 59200 46460 60000 46700
rect 0 46052 800 46292
rect 59200 45644 60000 45884
rect 0 45236 800 45476
rect 59200 44964 60000 45204
rect 0 44420 800 44660
rect 59200 44148 60000 44388
rect 0 43604 800 43844
rect 59200 43468 60000 43708
rect 0 42788 800 43028
rect 59200 42652 60000 42892
rect 0 41972 800 42212
rect 59200 41972 60000 42212
rect 0 41156 800 41396
rect 59200 41156 60000 41396
rect 0 40340 800 40580
rect 59200 40340 60000 40580
rect 0 39388 800 39628
rect 59200 39660 60000 39900
rect 0 38572 800 38812
rect 59200 38844 60000 39084
rect 59200 38164 60000 38404
rect 0 37756 800 37996
rect 59200 37348 60000 37588
rect 0 36940 800 37180
rect 59200 36532 60000 36772
rect 0 36124 800 36364
rect 59200 35852 60000 36092
rect 0 35308 800 35548
rect 59200 35036 60000 35276
rect 0 34492 800 34732
rect 59200 34356 60000 34596
rect 0 33676 800 33916
rect 59200 33540 60000 33780
rect 0 32724 800 32964
rect 59200 32860 60000 33100
rect 0 31908 800 32148
rect 59200 32044 60000 32284
rect 0 31092 800 31332
rect 59200 31228 60000 31468
rect 0 30276 800 30516
rect 59200 30548 60000 30788
rect 0 29460 800 29700
rect 59200 29732 60000 29972
rect 59200 29052 60000 29292
rect 0 28644 800 28884
rect 59200 28236 60000 28476
rect 0 27828 800 28068
rect 59200 27420 60000 27660
rect 0 27012 800 27252
rect 59200 26740 60000 26980
rect 0 26060 800 26300
rect 59200 25924 60000 26164
rect 0 25244 800 25484
rect 59200 25244 60000 25484
rect 0 24428 800 24668
rect 59200 24428 60000 24668
rect 0 23612 800 23852
rect 59200 23748 60000 23988
rect 0 22796 800 23036
rect 59200 22932 60000 23172
rect 0 21980 800 22220
rect 59200 22116 60000 22356
rect 0 21164 800 21404
rect 59200 21436 60000 21676
rect 0 20348 800 20588
rect 59200 20620 60000 20860
rect 59200 19940 60000 20180
rect 0 19396 800 19636
rect 59200 19124 60000 19364
rect 0 18580 800 18820
rect 59200 18308 60000 18548
rect 0 17764 800 18004
rect 59200 17628 60000 17868
rect 0 16948 800 17188
rect 59200 16812 60000 17052
rect 0 16132 800 16372
rect 59200 16132 60000 16372
rect 0 15316 800 15556
rect 59200 15316 60000 15556
rect 0 14500 800 14740
rect 59200 14636 60000 14876
rect 0 13684 800 13924
rect 59200 13820 60000 14060
rect 0 12732 800 12972
rect 59200 13004 60000 13244
rect 59200 12324 60000 12564
rect 0 11916 800 12156
rect 59200 11508 60000 11748
rect 0 11100 800 11340
rect 59200 10828 60000 11068
rect 0 10284 800 10524
rect 59200 10012 60000 10252
rect 0 9468 800 9708
rect 59200 9196 60000 9436
rect 0 8652 800 8892
rect 59200 8516 60000 8756
rect 0 7836 800 8076
rect 59200 7700 60000 7940
rect 0 7020 800 7260
rect 59200 7020 60000 7260
rect 0 6068 800 6308
rect 59200 6204 60000 6444
rect 0 5252 800 5492
rect 59200 5524 60000 5764
rect 0 4436 800 4676
rect 59200 4708 60000 4948
rect 0 3620 800 3860
rect 59200 3892 60000 4132
rect 59200 3212 60000 3452
rect 0 2804 800 3044
rect 59200 2396 60000 2636
rect 0 1988 800 2228
rect 59200 1716 60000 1956
rect 0 1172 800 1412
rect 59200 900 60000 1140
rect 0 356 800 596
rect 59200 220 60000 460
<< obsm3 >>
rect 880 59300 59120 59533
rect 800 58884 59200 59300
rect 880 58484 59120 58884
rect 800 58204 59200 58484
rect 800 58068 59120 58204
rect 880 57804 59120 58068
rect 880 57668 59200 57804
rect 800 57388 59200 57668
rect 800 57252 59120 57388
rect 880 56988 59120 57252
rect 880 56852 59200 56988
rect 800 56708 59200 56852
rect 800 56436 59120 56708
rect 880 56308 59120 56436
rect 880 56036 59200 56308
rect 800 55892 59200 56036
rect 800 55620 59120 55892
rect 880 55492 59120 55620
rect 880 55220 59200 55492
rect 800 55076 59200 55220
rect 800 54804 59120 55076
rect 880 54676 59120 54804
rect 880 54404 59200 54676
rect 800 54396 59200 54404
rect 800 53996 59120 54396
rect 800 53988 59200 53996
rect 880 53588 59200 53988
rect 800 53580 59200 53588
rect 800 53180 59120 53580
rect 800 53036 59200 53180
rect 880 52900 59200 53036
rect 880 52636 59120 52900
rect 800 52500 59120 52636
rect 800 52220 59200 52500
rect 880 52084 59200 52220
rect 880 51820 59120 52084
rect 800 51684 59120 51820
rect 800 51404 59200 51684
rect 880 51004 59120 51404
rect 800 50588 59200 51004
rect 880 50188 59120 50588
rect 800 49772 59200 50188
rect 880 49372 59120 49772
rect 800 49092 59200 49372
rect 800 48956 59120 49092
rect 880 48692 59120 48956
rect 880 48556 59200 48692
rect 800 48276 59200 48556
rect 800 48140 59120 48276
rect 880 47876 59120 48140
rect 880 47740 59200 47876
rect 800 47596 59200 47740
rect 800 47324 59120 47596
rect 880 47196 59120 47324
rect 880 46924 59200 47196
rect 800 46780 59200 46924
rect 800 46380 59120 46780
rect 800 46372 59200 46380
rect 880 45972 59200 46372
rect 800 45964 59200 45972
rect 800 45564 59120 45964
rect 800 45556 59200 45564
rect 880 45284 59200 45556
rect 880 45156 59120 45284
rect 800 44884 59120 45156
rect 800 44740 59200 44884
rect 880 44468 59200 44740
rect 880 44340 59120 44468
rect 800 44068 59120 44340
rect 800 43924 59200 44068
rect 880 43788 59200 43924
rect 880 43524 59120 43788
rect 800 43388 59120 43524
rect 800 43108 59200 43388
rect 880 42972 59200 43108
rect 880 42708 59120 42972
rect 800 42572 59120 42708
rect 800 42292 59200 42572
rect 880 41892 59120 42292
rect 800 41476 59200 41892
rect 880 41076 59120 41476
rect 800 40660 59200 41076
rect 880 40260 59120 40660
rect 800 39980 59200 40260
rect 800 39708 59120 39980
rect 880 39580 59120 39708
rect 880 39308 59200 39580
rect 800 39164 59200 39308
rect 800 38892 59120 39164
rect 880 38764 59120 38892
rect 880 38492 59200 38764
rect 800 38484 59200 38492
rect 800 38084 59120 38484
rect 800 38076 59200 38084
rect 880 37676 59200 38076
rect 800 37668 59200 37676
rect 800 37268 59120 37668
rect 800 37260 59200 37268
rect 880 36860 59200 37260
rect 800 36852 59200 36860
rect 800 36452 59120 36852
rect 800 36444 59200 36452
rect 880 36172 59200 36444
rect 880 36044 59120 36172
rect 800 35772 59120 36044
rect 800 35628 59200 35772
rect 880 35356 59200 35628
rect 880 35228 59120 35356
rect 800 34956 59120 35228
rect 800 34812 59200 34956
rect 880 34676 59200 34812
rect 880 34412 59120 34676
rect 800 34276 59120 34412
rect 800 33996 59200 34276
rect 880 33860 59200 33996
rect 880 33596 59120 33860
rect 800 33460 59120 33596
rect 800 33180 59200 33460
rect 800 33044 59120 33180
rect 880 32780 59120 33044
rect 880 32644 59200 32780
rect 800 32364 59200 32644
rect 800 32228 59120 32364
rect 880 31964 59120 32228
rect 880 31828 59200 31964
rect 800 31548 59200 31828
rect 800 31412 59120 31548
rect 880 31148 59120 31412
rect 880 31012 59200 31148
rect 800 30868 59200 31012
rect 800 30596 59120 30868
rect 880 30468 59120 30596
rect 880 30196 59200 30468
rect 800 30052 59200 30196
rect 800 29780 59120 30052
rect 880 29652 59120 29780
rect 880 29380 59200 29652
rect 800 29372 59200 29380
rect 800 28972 59120 29372
rect 800 28964 59200 28972
rect 880 28564 59200 28964
rect 800 28556 59200 28564
rect 800 28156 59120 28556
rect 800 28148 59200 28156
rect 880 27748 59200 28148
rect 800 27740 59200 27748
rect 800 27340 59120 27740
rect 800 27332 59200 27340
rect 880 27060 59200 27332
rect 880 26932 59120 27060
rect 800 26660 59120 26932
rect 800 26380 59200 26660
rect 880 26244 59200 26380
rect 880 25980 59120 26244
rect 800 25844 59120 25980
rect 800 25564 59200 25844
rect 880 25164 59120 25564
rect 800 24748 59200 25164
rect 880 24348 59120 24748
rect 800 24068 59200 24348
rect 800 23932 59120 24068
rect 880 23668 59120 23932
rect 880 23532 59200 23668
rect 800 23252 59200 23532
rect 800 23116 59120 23252
rect 880 22852 59120 23116
rect 880 22716 59200 22852
rect 800 22436 59200 22716
rect 800 22300 59120 22436
rect 880 22036 59120 22300
rect 880 21900 59200 22036
rect 800 21756 59200 21900
rect 800 21484 59120 21756
rect 880 21356 59120 21484
rect 880 21084 59200 21356
rect 800 20940 59200 21084
rect 800 20668 59120 20940
rect 880 20540 59120 20668
rect 880 20268 59200 20540
rect 800 20260 59200 20268
rect 800 19860 59120 20260
rect 800 19716 59200 19860
rect 880 19444 59200 19716
rect 880 19316 59120 19444
rect 800 19044 59120 19316
rect 800 18900 59200 19044
rect 880 18628 59200 18900
rect 880 18500 59120 18628
rect 800 18228 59120 18500
rect 800 18084 59200 18228
rect 880 17948 59200 18084
rect 880 17684 59120 17948
rect 800 17548 59120 17684
rect 800 17268 59200 17548
rect 880 17132 59200 17268
rect 880 16868 59120 17132
rect 800 16732 59120 16868
rect 800 16452 59200 16732
rect 880 16052 59120 16452
rect 800 15636 59200 16052
rect 880 15236 59120 15636
rect 800 14956 59200 15236
rect 800 14820 59120 14956
rect 880 14556 59120 14820
rect 880 14420 59200 14556
rect 800 14140 59200 14420
rect 800 14004 59120 14140
rect 880 13740 59120 14004
rect 880 13604 59200 13740
rect 800 13324 59200 13604
rect 800 13052 59120 13324
rect 880 12924 59120 13052
rect 880 12652 59200 12924
rect 800 12644 59200 12652
rect 800 12244 59120 12644
rect 800 12236 59200 12244
rect 880 11836 59200 12236
rect 800 11828 59200 11836
rect 800 11428 59120 11828
rect 800 11420 59200 11428
rect 880 11148 59200 11420
rect 880 11020 59120 11148
rect 800 10748 59120 11020
rect 800 10604 59200 10748
rect 880 10332 59200 10604
rect 880 10204 59120 10332
rect 800 9932 59120 10204
rect 800 9788 59200 9932
rect 880 9516 59200 9788
rect 880 9388 59120 9516
rect 800 9116 59120 9388
rect 800 8972 59200 9116
rect 880 8836 59200 8972
rect 880 8572 59120 8836
rect 800 8436 59120 8572
rect 800 8156 59200 8436
rect 880 8020 59200 8156
rect 880 7756 59120 8020
rect 800 7620 59120 7756
rect 800 7340 59200 7620
rect 880 6940 59120 7340
rect 800 6524 59200 6940
rect 800 6388 59120 6524
rect 880 6124 59120 6388
rect 880 5988 59200 6124
rect 800 5844 59200 5988
rect 800 5572 59120 5844
rect 880 5444 59120 5572
rect 880 5172 59200 5444
rect 800 5028 59200 5172
rect 800 4756 59120 5028
rect 880 4628 59120 4756
rect 880 4356 59200 4628
rect 800 4212 59200 4356
rect 800 3940 59120 4212
rect 880 3812 59120 3940
rect 880 3540 59200 3812
rect 800 3532 59200 3540
rect 800 3132 59120 3532
rect 800 3124 59200 3132
rect 880 2724 59200 3124
rect 800 2716 59200 2724
rect 800 2316 59120 2716
rect 800 2308 59200 2316
rect 880 2036 59200 2308
rect 880 1908 59120 2036
rect 800 1636 59120 1908
rect 800 1492 59200 1636
rect 880 1220 59200 1492
rect 880 1092 59120 1220
rect 800 820 59120 1092
rect 800 676 59200 820
rect 880 540 59200 676
rect 880 511 59120 540
<< metal4 >>
rect 4208 496 4528 57712
rect 19568 496 19888 57712
rect 34928 496 35248 57712
rect 50288 496 50608 57712
<< obsm4 >>
rect 12571 1259 19488 56677
rect 19968 1259 34848 56677
rect 35328 1259 45757 56677
<< labels >>
rlabel metal2 s 542 59200 654 60000 6 active
port 1 nsew signal input
rlabel metal2 s 2750 59200 2862 60000 6 io_in[0]
port 2 nsew signal input
rlabel metal2 s 14066 59200 14178 60000 6 io_in[10]
port 3 nsew signal input
rlabel metal2 s 15170 59200 15282 60000 6 io_in[11]
port 4 nsew signal input
rlabel metal2 s 16366 59200 16478 60000 6 io_in[12]
port 5 nsew signal input
rlabel metal2 s 17470 59200 17582 60000 6 io_in[13]
port 6 nsew signal input
rlabel metal2 s 18574 59200 18686 60000 6 io_in[14]
port 7 nsew signal input
rlabel metal2 s 19770 59200 19882 60000 6 io_in[15]
port 8 nsew signal input
rlabel metal2 s 20874 59200 20986 60000 6 io_in[16]
port 9 nsew signal input
rlabel metal2 s 21978 59200 22090 60000 6 io_in[17]
port 10 nsew signal input
rlabel metal2 s 23174 59200 23286 60000 6 io_in[18]
port 11 nsew signal input
rlabel metal2 s 24278 59200 24390 60000 6 io_in[19]
port 12 nsew signal input
rlabel metal2 s 3854 59200 3966 60000 6 io_in[1]
port 13 nsew signal input
rlabel metal2 s 25382 59200 25494 60000 6 io_in[20]
port 14 nsew signal input
rlabel metal2 s 26486 59200 26598 60000 6 io_in[21]
port 15 nsew signal input
rlabel metal2 s 27682 59200 27794 60000 6 io_in[22]
port 16 nsew signal input
rlabel metal2 s 28786 59200 28898 60000 6 io_in[23]
port 17 nsew signal input
rlabel metal2 s 29890 59200 30002 60000 6 io_in[24]
port 18 nsew signal input
rlabel metal2 s 31086 59200 31198 60000 6 io_in[25]
port 19 nsew signal input
rlabel metal2 s 32190 59200 32302 60000 6 io_in[26]
port 20 nsew signal input
rlabel metal2 s 33294 59200 33406 60000 6 io_in[27]
port 21 nsew signal input
rlabel metal2 s 34490 59200 34602 60000 6 io_in[28]
port 22 nsew signal input
rlabel metal2 s 35594 59200 35706 60000 6 io_in[29]
port 23 nsew signal input
rlabel metal2 s 5050 59200 5162 60000 6 io_in[2]
port 24 nsew signal input
rlabel metal2 s 36698 59200 36810 60000 6 io_in[30]
port 25 nsew signal input
rlabel metal2 s 37802 59200 37914 60000 6 io_in[31]
port 26 nsew signal input
rlabel metal2 s 38998 59200 39110 60000 6 io_in[32]
port 27 nsew signal input
rlabel metal2 s 40102 59200 40214 60000 6 io_in[33]
port 28 nsew signal input
rlabel metal2 s 41206 59200 41318 60000 6 io_in[34]
port 29 nsew signal input
rlabel metal2 s 42402 59200 42514 60000 6 io_in[35]
port 30 nsew signal input
rlabel metal2 s 43506 59200 43618 60000 6 io_in[36]
port 31 nsew signal input
rlabel metal2 s 44610 59200 44722 60000 6 io_in[37]
port 32 nsew signal input
rlabel metal2 s 6154 59200 6266 60000 6 io_in[3]
port 33 nsew signal input
rlabel metal2 s 7258 59200 7370 60000 6 io_in[4]
port 34 nsew signal input
rlabel metal2 s 8454 59200 8566 60000 6 io_in[5]
port 35 nsew signal input
rlabel metal2 s 9558 59200 9670 60000 6 io_in[6]
port 36 nsew signal input
rlabel metal2 s 10662 59200 10774 60000 6 io_in[7]
port 37 nsew signal input
rlabel metal2 s 11858 59200 11970 60000 6 io_in[8]
port 38 nsew signal input
rlabel metal2 s 12962 59200 13074 60000 6 io_in[9]
port 39 nsew signal input
rlabel metal3 s 59200 24428 60000 24668 6 io_oeb[0]
port 40 nsew signal output
rlabel metal3 s 59200 32044 60000 32284 6 io_oeb[10]
port 41 nsew signal output
rlabel metal3 s 59200 32860 60000 33100 6 io_oeb[11]
port 42 nsew signal output
rlabel metal3 s 59200 33540 60000 33780 6 io_oeb[12]
port 43 nsew signal output
rlabel metal3 s 59200 34356 60000 34596 6 io_oeb[13]
port 44 nsew signal output
rlabel metal3 s 59200 35036 60000 35276 6 io_oeb[14]
port 45 nsew signal output
rlabel metal3 s 59200 35852 60000 36092 6 io_oeb[15]
port 46 nsew signal output
rlabel metal3 s 59200 36532 60000 36772 6 io_oeb[16]
port 47 nsew signal output
rlabel metal3 s 59200 37348 60000 37588 6 io_oeb[17]
port 48 nsew signal output
rlabel metal3 s 59200 38164 60000 38404 6 io_oeb[18]
port 49 nsew signal output
rlabel metal3 s 59200 38844 60000 39084 6 io_oeb[19]
port 50 nsew signal output
rlabel metal3 s 59200 25244 60000 25484 6 io_oeb[1]
port 51 nsew signal output
rlabel metal3 s 59200 39660 60000 39900 6 io_oeb[20]
port 52 nsew signal output
rlabel metal3 s 59200 40340 60000 40580 6 io_oeb[21]
port 53 nsew signal output
rlabel metal3 s 59200 41156 60000 41396 6 io_oeb[22]
port 54 nsew signal output
rlabel metal3 s 59200 41972 60000 42212 6 io_oeb[23]
port 55 nsew signal output
rlabel metal3 s 59200 42652 60000 42892 6 io_oeb[24]
port 56 nsew signal output
rlabel metal3 s 59200 43468 60000 43708 6 io_oeb[25]
port 57 nsew signal output
rlabel metal3 s 59200 44148 60000 44388 6 io_oeb[26]
port 58 nsew signal output
rlabel metal3 s 59200 44964 60000 45204 6 io_oeb[27]
port 59 nsew signal output
rlabel metal3 s 59200 45644 60000 45884 6 io_oeb[28]
port 60 nsew signal output
rlabel metal3 s 59200 46460 60000 46700 6 io_oeb[29]
port 61 nsew signal output
rlabel metal3 s 59200 25924 60000 26164 6 io_oeb[2]
port 62 nsew signal output
rlabel metal3 s 59200 47276 60000 47516 6 io_oeb[30]
port 63 nsew signal output
rlabel metal3 s 59200 47956 60000 48196 6 io_oeb[31]
port 64 nsew signal output
rlabel metal3 s 59200 48772 60000 49012 6 io_oeb[32]
port 65 nsew signal output
rlabel metal3 s 59200 49452 60000 49692 6 io_oeb[33]
port 66 nsew signal output
rlabel metal3 s 59200 50268 60000 50508 6 io_oeb[34]
port 67 nsew signal output
rlabel metal3 s 59200 51084 60000 51324 6 io_oeb[35]
port 68 nsew signal output
rlabel metal3 s 59200 51764 60000 52004 6 io_oeb[36]
port 69 nsew signal output
rlabel metal3 s 59200 52580 60000 52820 6 io_oeb[37]
port 70 nsew signal output
rlabel metal3 s 59200 26740 60000 26980 6 io_oeb[3]
port 71 nsew signal output
rlabel metal3 s 59200 27420 60000 27660 6 io_oeb[4]
port 72 nsew signal output
rlabel metal3 s 59200 28236 60000 28476 6 io_oeb[5]
port 73 nsew signal output
rlabel metal3 s 59200 29052 60000 29292 6 io_oeb[6]
port 74 nsew signal output
rlabel metal3 s 59200 29732 60000 29972 6 io_oeb[7]
port 75 nsew signal output
rlabel metal3 s 59200 30548 60000 30788 6 io_oeb[8]
port 76 nsew signal output
rlabel metal3 s 59200 31228 60000 31468 6 io_oeb[9]
port 77 nsew signal output
rlabel metal2 s 45806 59200 45918 60000 6 io_out[0]
port 78 nsew signal output
rlabel metal2 s 11122 0 11234 800 6 io_out[10]
port 79 nsew signal output
rlabel metal3 s 59200 54076 60000 54316 6 io_out[11]
port 80 nsew signal output
rlabel metal2 s 18666 0 18778 800 6 io_out[12]
port 81 nsew signal output
rlabel metal2 s 26118 0 26230 800 6 io_out[13]
port 82 nsew signal output
rlabel metal2 s 33662 0 33774 800 6 io_out[14]
port 83 nsew signal output
rlabel metal3 s 0 56116 800 56356 6 io_out[15]
port 84 nsew signal output
rlabel metal3 s 59200 54756 60000 54996 6 io_out[16]
port 85 nsew signal output
rlabel metal2 s 41114 0 41226 800 6 io_out[17]
port 86 nsew signal output
rlabel metal2 s 51418 59200 51530 60000 6 io_out[18]
port 87 nsew signal output
rlabel metal3 s 59200 55572 60000 55812 6 io_out[19]
port 88 nsew signal output
rlabel metal2 s 46910 59200 47022 60000 6 io_out[1]
port 89 nsew signal output
rlabel metal2 s 48658 0 48770 800 6 io_out[20]
port 90 nsew signal output
rlabel metal2 s 52522 59200 52634 60000 6 io_out[21]
port 91 nsew signal output
rlabel metal2 s 53718 59200 53830 60000 6 io_out[22]
port 92 nsew signal output
rlabel metal2 s 54822 59200 54934 60000 6 io_out[23]
port 93 nsew signal output
rlabel metal3 s 0 56932 800 57172 6 io_out[24]
port 94 nsew signal output
rlabel metal3 s 59200 56388 60000 56628 6 io_out[25]
port 95 nsew signal output
rlabel metal2 s 55926 59200 56038 60000 6 io_out[26]
port 96 nsew signal output
rlabel metal3 s 59200 57068 60000 57308 6 io_out[27]
port 97 nsew signal output
rlabel metal3 s 0 57748 800 57988 6 io_out[28]
port 98 nsew signal output
rlabel metal3 s 59200 57884 60000 58124 6 io_out[29]
port 99 nsew signal output
rlabel metal2 s 48014 59200 48126 60000 6 io_out[2]
port 100 nsew signal output
rlabel metal2 s 56110 0 56222 800 6 io_out[30]
port 101 nsew signal output
rlabel metal2 s 57122 59200 57234 60000 6 io_out[31]
port 102 nsew signal output
rlabel metal2 s 58226 59200 58338 60000 6 io_out[32]
port 103 nsew signal output
rlabel metal3 s 0 58564 800 58804 6 io_out[33]
port 104 nsew signal output
rlabel metal3 s 59200 58564 60000 58804 6 io_out[34]
port 105 nsew signal output
rlabel metal3 s 0 59380 800 59620 6 io_out[35]
port 106 nsew signal output
rlabel metal3 s 59200 59380 60000 59620 6 io_out[36]
port 107 nsew signal output
rlabel metal2 s 59330 59200 59442 60000 6 io_out[37]
port 108 nsew signal output
rlabel metal2 s 3670 0 3782 800 6 io_out[3]
port 109 nsew signal output
rlabel metal3 s 0 53668 800 53908 6 io_out[4]
port 110 nsew signal output
rlabel metal3 s 59200 53260 60000 53500 6 io_out[5]
port 111 nsew signal output
rlabel metal3 s 0 54484 800 54724 6 io_out[6]
port 112 nsew signal output
rlabel metal2 s 49118 59200 49230 60000 6 io_out[7]
port 113 nsew signal output
rlabel metal2 s 50314 59200 50426 60000 6 io_out[8]
port 114 nsew signal output
rlabel metal3 s 0 55300 800 55540 6 io_out[9]
port 115 nsew signal output
rlabel metal3 s 0 356 800 596 6 la1_data_in[0]
port 116 nsew signal input
rlabel metal3 s 0 8652 800 8892 6 la1_data_in[10]
port 117 nsew signal input
rlabel metal3 s 0 9468 800 9708 6 la1_data_in[11]
port 118 nsew signal input
rlabel metal3 s 0 10284 800 10524 6 la1_data_in[12]
port 119 nsew signal input
rlabel metal3 s 0 11100 800 11340 6 la1_data_in[13]
port 120 nsew signal input
rlabel metal3 s 0 11916 800 12156 6 la1_data_in[14]
port 121 nsew signal input
rlabel metal3 s 0 12732 800 12972 6 la1_data_in[15]
port 122 nsew signal input
rlabel metal3 s 0 13684 800 13924 6 la1_data_in[16]
port 123 nsew signal input
rlabel metal3 s 0 14500 800 14740 6 la1_data_in[17]
port 124 nsew signal input
rlabel metal3 s 0 15316 800 15556 6 la1_data_in[18]
port 125 nsew signal input
rlabel metal3 s 0 16132 800 16372 6 la1_data_in[19]
port 126 nsew signal input
rlabel metal3 s 0 1172 800 1412 6 la1_data_in[1]
port 127 nsew signal input
rlabel metal3 s 0 16948 800 17188 6 la1_data_in[20]
port 128 nsew signal input
rlabel metal3 s 0 17764 800 18004 6 la1_data_in[21]
port 129 nsew signal input
rlabel metal3 s 0 18580 800 18820 6 la1_data_in[22]
port 130 nsew signal input
rlabel metal3 s 0 19396 800 19636 6 la1_data_in[23]
port 131 nsew signal input
rlabel metal3 s 0 20348 800 20588 6 la1_data_in[24]
port 132 nsew signal input
rlabel metal3 s 0 21164 800 21404 6 la1_data_in[25]
port 133 nsew signal input
rlabel metal3 s 0 21980 800 22220 6 la1_data_in[26]
port 134 nsew signal input
rlabel metal3 s 0 22796 800 23036 6 la1_data_in[27]
port 135 nsew signal input
rlabel metal3 s 0 23612 800 23852 6 la1_data_in[28]
port 136 nsew signal input
rlabel metal3 s 0 24428 800 24668 6 la1_data_in[29]
port 137 nsew signal input
rlabel metal3 s 0 1988 800 2228 6 la1_data_in[2]
port 138 nsew signal input
rlabel metal3 s 0 25244 800 25484 6 la1_data_in[30]
port 139 nsew signal input
rlabel metal3 s 0 26060 800 26300 6 la1_data_in[31]
port 140 nsew signal input
rlabel metal3 s 0 2804 800 3044 6 la1_data_in[3]
port 141 nsew signal input
rlabel metal3 s 0 3620 800 3860 6 la1_data_in[4]
port 142 nsew signal input
rlabel metal3 s 0 4436 800 4676 6 la1_data_in[5]
port 143 nsew signal input
rlabel metal3 s 0 5252 800 5492 6 la1_data_in[6]
port 144 nsew signal input
rlabel metal3 s 0 6068 800 6308 6 la1_data_in[7]
port 145 nsew signal input
rlabel metal3 s 0 7020 800 7260 6 la1_data_in[8]
port 146 nsew signal input
rlabel metal3 s 0 7836 800 8076 6 la1_data_in[9]
port 147 nsew signal input
rlabel metal3 s 0 27012 800 27252 6 la1_data_out[0]
port 148 nsew signal output
rlabel metal3 s 0 35308 800 35548 6 la1_data_out[10]
port 149 nsew signal output
rlabel metal3 s 0 36124 800 36364 6 la1_data_out[11]
port 150 nsew signal output
rlabel metal3 s 0 36940 800 37180 6 la1_data_out[12]
port 151 nsew signal output
rlabel metal3 s 0 37756 800 37996 6 la1_data_out[13]
port 152 nsew signal output
rlabel metal3 s 0 38572 800 38812 6 la1_data_out[14]
port 153 nsew signal output
rlabel metal3 s 0 39388 800 39628 6 la1_data_out[15]
port 154 nsew signal output
rlabel metal3 s 0 40340 800 40580 6 la1_data_out[16]
port 155 nsew signal output
rlabel metal3 s 0 41156 800 41396 6 la1_data_out[17]
port 156 nsew signal output
rlabel metal3 s 0 41972 800 42212 6 la1_data_out[18]
port 157 nsew signal output
rlabel metal3 s 0 42788 800 43028 6 la1_data_out[19]
port 158 nsew signal output
rlabel metal3 s 0 27828 800 28068 6 la1_data_out[1]
port 159 nsew signal output
rlabel metal3 s 0 43604 800 43844 6 la1_data_out[20]
port 160 nsew signal output
rlabel metal3 s 0 44420 800 44660 6 la1_data_out[21]
port 161 nsew signal output
rlabel metal3 s 0 45236 800 45476 6 la1_data_out[22]
port 162 nsew signal output
rlabel metal3 s 0 46052 800 46292 6 la1_data_out[23]
port 163 nsew signal output
rlabel metal3 s 0 47004 800 47244 6 la1_data_out[24]
port 164 nsew signal output
rlabel metal3 s 0 47820 800 48060 6 la1_data_out[25]
port 165 nsew signal output
rlabel metal3 s 0 48636 800 48876 6 la1_data_out[26]
port 166 nsew signal output
rlabel metal3 s 0 49452 800 49692 6 la1_data_out[27]
port 167 nsew signal output
rlabel metal3 s 0 50268 800 50508 6 la1_data_out[28]
port 168 nsew signal output
rlabel metal3 s 0 51084 800 51324 6 la1_data_out[29]
port 169 nsew signal output
rlabel metal3 s 0 28644 800 28884 6 la1_data_out[2]
port 170 nsew signal output
rlabel metal3 s 0 51900 800 52140 6 la1_data_out[30]
port 171 nsew signal output
rlabel metal3 s 0 52716 800 52956 6 la1_data_out[31]
port 172 nsew signal output
rlabel metal3 s 0 29460 800 29700 6 la1_data_out[3]
port 173 nsew signal output
rlabel metal3 s 0 30276 800 30516 6 la1_data_out[4]
port 174 nsew signal output
rlabel metal3 s 0 31092 800 31332 6 la1_data_out[5]
port 175 nsew signal output
rlabel metal3 s 0 31908 800 32148 6 la1_data_out[6]
port 176 nsew signal output
rlabel metal3 s 0 32724 800 32964 6 la1_data_out[7]
port 177 nsew signal output
rlabel metal3 s 0 33676 800 33916 6 la1_data_out[8]
port 178 nsew signal output
rlabel metal3 s 0 34492 800 34732 6 la1_data_out[9]
port 179 nsew signal output
rlabel metal3 s 59200 220 60000 460 6 la1_oenb[0]
port 180 nsew signal input
rlabel metal3 s 59200 7700 60000 7940 6 la1_oenb[10]
port 181 nsew signal input
rlabel metal3 s 59200 8516 60000 8756 6 la1_oenb[11]
port 182 nsew signal input
rlabel metal3 s 59200 9196 60000 9436 6 la1_oenb[12]
port 183 nsew signal input
rlabel metal3 s 59200 10012 60000 10252 6 la1_oenb[13]
port 184 nsew signal input
rlabel metal3 s 59200 10828 60000 11068 6 la1_oenb[14]
port 185 nsew signal input
rlabel metal3 s 59200 11508 60000 11748 6 la1_oenb[15]
port 186 nsew signal input
rlabel metal3 s 59200 12324 60000 12564 6 la1_oenb[16]
port 187 nsew signal input
rlabel metal3 s 59200 13004 60000 13244 6 la1_oenb[17]
port 188 nsew signal input
rlabel metal3 s 59200 13820 60000 14060 6 la1_oenb[18]
port 189 nsew signal input
rlabel metal3 s 59200 14636 60000 14876 6 la1_oenb[19]
port 190 nsew signal input
rlabel metal3 s 59200 900 60000 1140 6 la1_oenb[1]
port 191 nsew signal input
rlabel metal3 s 59200 15316 60000 15556 6 la1_oenb[20]
port 192 nsew signal input
rlabel metal3 s 59200 16132 60000 16372 6 la1_oenb[21]
port 193 nsew signal input
rlabel metal3 s 59200 16812 60000 17052 6 la1_oenb[22]
port 194 nsew signal input
rlabel metal3 s 59200 17628 60000 17868 6 la1_oenb[23]
port 195 nsew signal input
rlabel metal3 s 59200 18308 60000 18548 6 la1_oenb[24]
port 196 nsew signal input
rlabel metal3 s 59200 19124 60000 19364 6 la1_oenb[25]
port 197 nsew signal input
rlabel metal3 s 59200 19940 60000 20180 6 la1_oenb[26]
port 198 nsew signal input
rlabel metal3 s 59200 20620 60000 20860 6 la1_oenb[27]
port 199 nsew signal input
rlabel metal3 s 59200 21436 60000 21676 6 la1_oenb[28]
port 200 nsew signal input
rlabel metal3 s 59200 22116 60000 22356 6 la1_oenb[29]
port 201 nsew signal input
rlabel metal3 s 59200 1716 60000 1956 6 la1_oenb[2]
port 202 nsew signal input
rlabel metal3 s 59200 22932 60000 23172 6 la1_oenb[30]
port 203 nsew signal input
rlabel metal3 s 59200 23748 60000 23988 6 la1_oenb[31]
port 204 nsew signal input
rlabel metal3 s 59200 2396 60000 2636 6 la1_oenb[3]
port 205 nsew signal input
rlabel metal3 s 59200 3212 60000 3452 6 la1_oenb[4]
port 206 nsew signal input
rlabel metal3 s 59200 3892 60000 4132 6 la1_oenb[5]
port 207 nsew signal input
rlabel metal3 s 59200 4708 60000 4948 6 la1_oenb[6]
port 208 nsew signal input
rlabel metal3 s 59200 5524 60000 5764 6 la1_oenb[7]
port 209 nsew signal input
rlabel metal3 s 59200 6204 60000 6444 6 la1_oenb[8]
port 210 nsew signal input
rlabel metal3 s 59200 7020 60000 7260 6 la1_oenb[9]
port 211 nsew signal input
rlabel metal4 s 4208 496 4528 57712 6 vccd1
port 212 nsew power input
rlabel metal4 s 34928 496 35248 57712 6 vccd1
port 212 nsew power input
rlabel metal4 s 19568 496 19888 57712 6 vssd1
port 213 nsew ground input
rlabel metal4 s 50288 496 50608 57712 6 vssd1
port 213 nsew ground input
rlabel metal2 s 1646 59200 1758 60000 6 wb_clk_i
port 214 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 60000 60000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 12364314
string GDS_FILE /openlane/designs/wrapped-vgademo-on-fpga/runs/RUN_2022.03.20_07.43.13/results/finishing/wrapped_vgademo_on_fpga.magic.gds
string GDS_START 1090352
<< end >>

