* NGSPICE file created from wrapped_vgademo_on_fpga.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_8 abstract view
.subckt sky130_fd_sc_hd__ebufn_8 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_4 abstract view
.subckt sky130_fd_sc_hd__nor2b_4 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_2 abstract view
.subckt sky130_fd_sc_hd__o32ai_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_4 abstract view
.subckt sky130_fd_sc_hd__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

.subckt wrapped_vgademo_on_fpga active io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21]
+ io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29]
+ io_in[2] io_in[30] io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37]
+ io_in[3] io_in[4] io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10]
+ io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18]
+ io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25]
+ io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32]
+ io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5]
+ io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12]
+ io_out[13] io_out[14] io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1]
+ io_out[20] io_out[21] io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27]
+ io_out[28] io_out[29] io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34]
+ io_out[35] io_out[36] io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ io_out[8] io_out[9] la1_data_in[0] la1_data_in[10] la1_data_in[11] la1_data_in[12]
+ la1_data_in[13] la1_data_in[14] la1_data_in[15] la1_data_in[16] la1_data_in[17]
+ la1_data_in[18] la1_data_in[19] la1_data_in[1] la1_data_in[20] la1_data_in[21] la1_data_in[22]
+ la1_data_in[23] la1_data_in[24] la1_data_in[25] la1_data_in[26] la1_data_in[27]
+ la1_data_in[28] la1_data_in[29] la1_data_in[2] la1_data_in[30] la1_data_in[31] la1_data_in[3]
+ la1_data_in[4] la1_data_in[5] la1_data_in[6] la1_data_in[7] la1_data_in[8] la1_data_in[9]
+ la1_data_out[0] la1_data_out[10] la1_data_out[11] la1_data_out[12] la1_data_out[13]
+ la1_data_out[14] la1_data_out[15] la1_data_out[16] la1_data_out[17] la1_data_out[18]
+ la1_data_out[19] la1_data_out[1] la1_data_out[20] la1_data_out[21] la1_data_out[22]
+ la1_data_out[23] la1_data_out[24] la1_data_out[25] la1_data_out[26] la1_data_out[27]
+ la1_data_out[28] la1_data_out[29] la1_data_out[2] la1_data_out[30] la1_data_out[31]
+ la1_data_out[3] la1_data_out[4] la1_data_out[5] la1_data_out[6] la1_data_out[7]
+ la1_data_out[8] la1_data_out[9] la1_oenb[0] la1_oenb[10] la1_oenb[11] la1_oenb[12]
+ la1_oenb[13] la1_oenb[14] la1_oenb[15] la1_oenb[16] la1_oenb[17] la1_oenb[18] la1_oenb[19]
+ la1_oenb[1] la1_oenb[20] la1_oenb[21] la1_oenb[22] la1_oenb[23] la1_oenb[24] la1_oenb[25]
+ la1_oenb[26] la1_oenb[27] la1_oenb[28] la1_oenb[29] la1_oenb[2] la1_oenb[30] la1_oenb[31]
+ la1_oenb[3] la1_oenb[4] la1_oenb[5] la1_oenb[6] la1_oenb[7] la1_oenb[8] la1_oenb[9]
+ vccd1 vssd1 wb_clk_i
XFILLER_79_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7963_ _8056_/A _7963_/B vssd1 vssd1 vccd1 vccd1 _7964_/C sky130_fd_sc_hd__nor2_1
XFILLER_27_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6914_ _6914_/A _7017_/B vssd1 vssd1 vccd1 vccd1 _6916_/A sky130_fd_sc_hd__xnor2_2
X_7894_ _7834_/A _7894_/B vssd1 vssd1 vccd1 vccd1 _7981_/A sky130_fd_sc_hd__and2b_1
XFILLER_23_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6845_ _6963_/A _6845_/B vssd1 vssd1 vccd1 vccd1 _6976_/B sky130_fd_sc_hd__xnor2_2
X_6776_ _7118_/B _6780_/A vssd1 vssd1 vccd1 vccd1 _6863_/B sky130_fd_sc_hd__nor2_1
X_8515_ _8461_/S _8513_/A _8513_/Y _8514_/X vssd1 vssd1 vccd1 vccd1 _8519_/A sky130_fd_sc_hd__a22o_1
X_5727_ _5727_/A _5727_/B _5741_/A vssd1 vssd1 vccd1 vccd1 _5728_/C sky130_fd_sc_hd__and3_1
X_8446_ _8399_/A _8398_/B _8396_/X vssd1 vssd1 vccd1 vccd1 _8469_/A sky130_fd_sc_hd__a21o_1
X_5658_ _5764_/A _5764_/B vssd1 vssd1 vccd1 vccd1 _5787_/A sky130_fd_sc_hd__xnor2_1
X_8377_ _7934_/B _8460_/A _7999_/X vssd1 vssd1 vccd1 vccd1 _8384_/A sky130_fd_sc_hd__a21o_1
X_5589_ _5892_/A vssd1 vssd1 vccd1 vccd1 _5984_/C sky130_fd_sc_hd__clkbuf_2
X_4609_ _8646_/Q _8645_/Q _8648_/Q _8651_/Q vssd1 vssd1 vccd1 vccd1 _4611_/C sky130_fd_sc_hd__or4b_1
X_7328_ _7309_/A _6813_/B _7231_/B _7327_/X vssd1 vssd1 vccd1 vccd1 _7335_/A sky130_fd_sc_hd__a31o_1
XFILLER_104_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7259_ _7259_/A _7195_/B vssd1 vssd1 vccd1 vccd1 _7259_/X sky130_fd_sc_hd__or2b_1
XFILLER_89_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4960_ _4995_/A _4960_/B vssd1 vssd1 vccd1 vccd1 _4980_/C sky130_fd_sc_hd__nand2_1
XFILLER_17_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4891_ _5033_/A _4891_/B vssd1 vssd1 vccd1 vccd1 _5154_/A sky130_fd_sc_hd__or2_1
XFILLER_20_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6630_ _8749_/Q _6630_/B vssd1 vssd1 vccd1 vccd1 _6630_/X sky130_fd_sc_hd__and2b_1
X_6561_ _6555_/X _6560_/Y _7621_/A vssd1 vssd1 vccd1 vccd1 _8747_/D sky130_fd_sc_hd__o21ai_1
X_8300_ _8345_/A _8300_/B vssd1 vssd1 vccd1 vccd1 _8302_/C sky130_fd_sc_hd__and2b_1
X_5512_ _6378_/A _5512_/B vssd1 vssd1 vccd1 vccd1 _5681_/A sky130_fd_sc_hd__nor2_2
X_6492_ _8734_/Q _8733_/Q _6492_/C vssd1 vssd1 vccd1 vccd1 _6497_/C sky130_fd_sc_hd__and3_1
X_8231_ _8222_/A _8222_/B _8221_/A vssd1 vssd1 vccd1 vccd1 _8308_/A sky130_fd_sc_hd__o21ai_2
X_5443_ _6460_/A _5443_/B vssd1 vssd1 vccd1 vccd1 _5449_/A sky130_fd_sc_hd__and2_1
X_8818__35 vssd1 vssd1 vccd1 vccd1 _8818__35/HI _8913_/A sky130_fd_sc_hd__conb_1
X_8162_ _8182_/A _8514_/B vssd1 vssd1 vccd1 vccd1 _8163_/B sky130_fd_sc_hd__or2_1
X_5374_ _5377_/C _5374_/B vssd1 vssd1 vccd1 vccd1 _8691_/D sky130_fd_sc_hd__nor2_1
X_7113_ _7116_/B _7116_/A vssd1 vssd1 vccd1 vccd1 _7113_/X sky130_fd_sc_hd__and2b_1
X_8093_ _8330_/A _8348_/B vssd1 vssd1 vccd1 vccd1 _8420_/A sky130_fd_sc_hd__or2_2
XFILLER_86_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7044_ _7165_/A _7165_/B vssd1 vssd1 vccd1 vccd1 _7061_/A sky130_fd_sc_hd__xor2_1
XFILLER_101_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7946_ _7946_/A _8348_/B vssd1 vssd1 vccd1 vccd1 _8120_/A sky130_fd_sc_hd__nor2_1
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7877_ _8325_/A _8325_/B vssd1 vssd1 vccd1 vccd1 _7878_/C sky130_fd_sc_hd__nand2_1
XFILLER_11_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6828_ _6898_/A _6966_/B _6965_/A vssd1 vssd1 vccd1 vccd1 _6829_/B sky130_fd_sc_hd__or3b_1
XFILLER_50_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6759_ _6775_/A _6775_/B _6755_/X vssd1 vssd1 vccd1 vccd1 _6759_/X sky130_fd_sc_hd__a21o_1
XFILLER_10_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8429_ _8506_/B _8429_/B vssd1 vssd1 vccd1 vccd1 _8433_/A sky130_fd_sc_hd__xnor2_1
XFILLER_12_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5090_ _5108_/B _5156_/B vssd1 vssd1 vccd1 vccd1 _5099_/D sky130_fd_sc_hd__or2_1
XFILLER_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7800_ _8273_/A _8172_/A vssd1 vssd1 vccd1 vccd1 _7800_/Y sky130_fd_sc_hd__nand2_1
X_5992_ _6183_/A _6192_/B vssd1 vssd1 vccd1 vccd1 _5995_/A sky130_fd_sc_hd__nor2_1
X_8780_ _8783_/CLK _8780_/D vssd1 vssd1 vccd1 vccd1 _8780_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7731_ _8782_/Q _8658_/Q vssd1 vssd1 vccd1 vccd1 _7733_/A sky130_fd_sc_hd__and2b_1
X_4943_ _4956_/A _5153_/C vssd1 vssd1 vccd1 vccd1 _4966_/A sky130_fd_sc_hd__or2_1
X_7662_ _7662_/A _7662_/B vssd1 vssd1 vccd1 vccd1 _7662_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_20_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6613_ _8760_/Q _6613_/B vssd1 vssd1 vccd1 vccd1 _6613_/X sky130_fd_sc_hd__and2b_1
X_4874_ _4874_/A _4874_/B vssd1 vssd1 vccd1 vccd1 _5298_/B sky130_fd_sc_hd__nor2_1
X_7593_ _8779_/Q vssd1 vssd1 vccd1 vccd1 _8595_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_20_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6544_ _8764_/Q vssd1 vssd1 vccd1 vccd1 _7583_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6475_ _6475_/A vssd1 vssd1 vccd1 vccd1 _8728_/D sky130_fd_sc_hd__clkbuf_1
X_8214_ _8214_/A _8214_/B _8214_/C vssd1 vssd1 vccd1 vccd1 _8214_/Y sky130_fd_sc_hd__nor3_1
X_5426_ _6415_/B vssd1 vssd1 vccd1 vccd1 _6427_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_8145_ _8118_/B _8145_/B vssd1 vssd1 vccd1 vccd1 _8145_/X sky130_fd_sc_hd__and2b_1
X_5357_ _5359_/B _5389_/B _5357_/C vssd1 vssd1 vccd1 vccd1 _5358_/A sky130_fd_sc_hd__and3b_1
XFILLER_87_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8076_ _8181_/A _8181_/B vssd1 vssd1 vccd1 vccd1 _8078_/B sky130_fd_sc_hd__xor2_1
X_5288_ _5288_/A _5288_/B _5288_/C vssd1 vssd1 vccd1 vccd1 _5288_/X sky130_fd_sc_hd__or3_1
XINSDIODE2_4 _5251_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7027_ _7027_/A _6916_/A vssd1 vssd1 vccd1 vccd1 _7041_/A sky130_fd_sc_hd__or2b_1
XFILLER_101_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8978_ _8978_/A _4473_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[27] sky130_fd_sc_hd__ebufn_8
XFILLER_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7929_ _8018_/A _7929_/B vssd1 vssd1 vccd1 vccd1 _7930_/C sky130_fd_sc_hd__and2b_1
XFILLER_55_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4590_ _4590_/A vssd1 vssd1 vccd1 vccd1 _8936_/A sky130_fd_sc_hd__clkbuf_1
X_6260_ _6199_/B _6260_/B vssd1 vssd1 vccd1 vccd1 _6268_/B sky130_fd_sc_hd__and2b_1
X_6191_ _6092_/A _6200_/B _5827_/X vssd1 vssd1 vccd1 vccd1 _6259_/A sky130_fd_sc_hd__a21o_1
X_5211_ _5211_/A _5211_/B _5211_/C _5211_/D vssd1 vssd1 vccd1 vccd1 _5211_/X sky130_fd_sc_hd__or4_1
X_5142_ _5250_/C _5149_/C _5142_/C _5088_/A vssd1 vssd1 vccd1 vccd1 _5142_/Y sky130_fd_sc_hd__nor4b_1
XFILLER_96_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5073_ _5073_/A _5073_/B _5073_/C vssd1 vssd1 vccd1 vccd1 _5073_/X sky130_fd_sc_hd__or3_1
X_8901_ _8901_/A _4382_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[20] sky130_fd_sc_hd__ebufn_8
XFILLER_37_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5975_ _5975_/A _5975_/B vssd1 vssd1 vccd1 vccd1 _5975_/Y sky130_fd_sc_hd__nand2_1
X_8763_ _8763_/CLK _8763_/D vssd1 vssd1 vccd1 vccd1 _8763_/Q sky130_fd_sc_hd__dfxtp_1
X_7714_ _7761_/A _7714_/B vssd1 vssd1 vccd1 vccd1 _7764_/B sky130_fd_sc_hd__xnor2_1
X_4926_ _5082_/B _4926_/B vssd1 vssd1 vccd1 vccd1 _5076_/A sky130_fd_sc_hd__nor2_1
X_8694_ _8704_/CLK _8694_/D vssd1 vssd1 vccd1 vccd1 _8694_/Q sky130_fd_sc_hd__dfxtp_1
X_7645_ _7649_/A _8767_/Q vssd1 vssd1 vccd1 vccd1 _7652_/B sky130_fd_sc_hd__xnor2_1
XFILLER_20_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4857_ _5078_/B vssd1 vssd1 vccd1 vccd1 _5174_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7576_ _7585_/A _7576_/B _7583_/B vssd1 vssd1 vccd1 vccd1 _7576_/X sky130_fd_sc_hd__and3_1
X_4788_ _4788_/A vssd1 vssd1 vccd1 vccd1 _8665_/D sky130_fd_sc_hd__clkbuf_1
X_6527_ _6653_/A vssd1 vssd1 vccd1 vccd1 _7587_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6458_ _7619_/B _7619_/C vssd1 vssd1 vccd1 vccd1 _7622_/B sky130_fd_sc_hd__nor2_1
X_6389_ _6388_/B _6389_/B vssd1 vssd1 vccd1 vccd1 _6390_/D sky130_fd_sc_hd__and2b_1
X_5409_ _5409_/A _5409_/B _5409_/C vssd1 vssd1 vccd1 vccd1 _5410_/A sky130_fd_sc_hd__and3_1
XFILLER_102_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8128_ _8128_/A _8128_/B vssd1 vssd1 vccd1 vccd1 _8129_/B sky130_fd_sc_hd__or2_1
XFILLER_87_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8059_ _8059_/A _8059_/B vssd1 vssd1 vccd1 vccd1 _8147_/A sky130_fd_sc_hd__nand2_1
XFILLER_18_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5760_ _6071_/A _6197_/A _5760_/C _5760_/D vssd1 vssd1 vccd1 vccd1 _5810_/B sky130_fd_sc_hd__nand4_2
XFILLER_22_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5691_ _5891_/A _5645_/C _5704_/A _5704_/B vssd1 vssd1 vccd1 vccd1 _5693_/B sky130_fd_sc_hd__o22a_1
XFILLER_30_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4711_ _5264_/A vssd1 vssd1 vccd1 vccd1 _5182_/A sky130_fd_sc_hd__buf_2
X_7430_ _7430_/A _7430_/B vssd1 vssd1 vccd1 vccd1 _7442_/B sky130_fd_sc_hd__xnor2_2
X_4642_ _8638_/Q _4643_/C _4641_/Y vssd1 vssd1 vccd1 vccd1 _8638_/D sky130_fd_sc_hd__a21oi_1
XFILLER_30_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7361_ _7434_/A _7508_/A vssd1 vssd1 vccd1 vccd1 _7361_/X sky130_fd_sc_hd__or2_1
X_4573_ _4573_/A _4573_/B _4702_/A vssd1 vssd1 vccd1 vccd1 _4574_/D sky130_fd_sc_hd__and3_1
X_6312_ _6249_/A _6173_/A _6312_/S vssd1 vssd1 vccd1 vccd1 _6313_/B sky130_fd_sc_hd__mux2_1
X_7292_ _7290_/Y _7292_/B vssd1 vssd1 vccd1 vccd1 _7293_/B sky130_fd_sc_hd__and2b_1
X_6243_ _6243_/A vssd1 vssd1 vccd1 vccd1 _6243_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6174_ _6166_/A _6251_/B _6302_/B _6224_/A vssd1 vssd1 vccd1 vccd1 _6175_/B sky130_fd_sc_hd__o22a_1
X_5125_ _5066_/A _5221_/C _5123_/X _5124_/X _5050_/D vssd1 vssd1 vccd1 vccd1 _5127_/B
+ sky130_fd_sc_hd__o32a_1
X_5056_ _5255_/A _5051_/X _5055_/X vssd1 vssd1 vccd1 vccd1 _5056_/X sky130_fd_sc_hd__o21a_1
XFILLER_37_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5958_ _6128_/A _6128_/B vssd1 vssd1 vccd1 vccd1 _6370_/B sky130_fd_sc_hd__xor2_2
XFILLER_52_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8746_ _8753_/CLK _8746_/D vssd1 vssd1 vccd1 vccd1 _8746_/Q sky130_fd_sc_hd__dfxtp_1
X_4909_ _4784_/A _4883_/B _5040_/B vssd1 vssd1 vccd1 vccd1 _5190_/A sky130_fd_sc_hd__a21oi_2
X_5889_ _5889_/A _5889_/B vssd1 vssd1 vccd1 vccd1 _5975_/A sky130_fd_sc_hd__nand2_1
X_8677_ _8776_/CLK _8677_/D vssd1 vssd1 vccd1 vccd1 _8677_/Q sky130_fd_sc_hd__dfxtp_1
X_7628_ _8628_/A vssd1 vssd1 vccd1 vccd1 _8603_/A sky130_fd_sc_hd__clkbuf_2
X_7559_ _7557_/Y _7559_/B vssd1 vssd1 vccd1 vccd1 _7559_/X sky130_fd_sc_hd__and2b_1
XFILLER_20_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8793__10 vssd1 vssd1 vccd1 vccd1 _8793__10/HI _8888_/A sky130_fd_sc_hd__conb_1
XFILLER_54_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6930_ _7030_/A _7302_/A vssd1 vssd1 vccd1 vccd1 _6943_/A sky130_fd_sc_hd__nor2_2
XFILLER_35_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6861_ _6861_/A _6861_/B vssd1 vssd1 vccd1 vccd1 _6879_/A sky130_fd_sc_hd__nor2_1
X_8600_ _8600_/A _8600_/B vssd1 vssd1 vccd1 vccd1 _8602_/A sky130_fd_sc_hd__nor2_1
X_5812_ _6071_/A _6197_/A _5760_/D _5811_/X vssd1 vssd1 vccd1 vccd1 _5847_/A sky130_fd_sc_hd__a31o_1
XFILLER_62_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6792_ _6836_/A _6792_/B vssd1 vssd1 vccd1 vccd1 _7262_/B sky130_fd_sc_hd__nand2_2
X_8531_ _8531_/A _8531_/B vssd1 vssd1 vccd1 vccd1 _8532_/B sky130_fd_sc_hd__xnor2_1
X_5743_ _5743_/A _5743_/B vssd1 vssd1 vccd1 vccd1 _5744_/C sky130_fd_sc_hd__xor2_1
X_8462_ _8513_/A _8513_/B vssd1 vssd1 vccd1 vccd1 _8465_/A sky130_fd_sc_hd__xnor2_1
X_5674_ _5679_/A _5715_/A _5674_/C vssd1 vssd1 vccd1 vccd1 _5676_/A sky130_fd_sc_hd__or3_1
XFILLER_30_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8393_ _8393_/A _8457_/B vssd1 vssd1 vccd1 vccd1 _8394_/C sky130_fd_sc_hd__xnor2_1
X_7413_ _7176_/A _7080_/C _7006_/X vssd1 vssd1 vccd1 vccd1 _7413_/Y sky130_fd_sc_hd__a21oi_1
X_4625_ _4625_/A vssd1 vssd1 vccd1 vccd1 _8633_/D sky130_fd_sc_hd__clkbuf_1
X_4556_ _8654_/Q vssd1 vssd1 vccd1 vccd1 _4733_/C sky130_fd_sc_hd__clkbuf_2
X_7344_ _7344_/A _7344_/B vssd1 vssd1 vccd1 vccd1 _7345_/B sky130_fd_sc_hd__xnor2_1
X_4487_ _4489_/A vssd1 vssd1 vccd1 vccd1 _4487_/Y sky130_fd_sc_hd__inv_2
XFILLER_89_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7275_ _6792_/B _7501_/A _7177_/B _7405_/A vssd1 vssd1 vccd1 vccd1 _7276_/C sky130_fd_sc_hd__a22o_1
XFILLER_103_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6226_ _6175_/A _6175_/B _6251_/B _6249_/A vssd1 vssd1 vccd1 vccd1 _6233_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_103_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6157_ _6157_/A _6113_/B vssd1 vssd1 vccd1 vccd1 _6158_/B sky130_fd_sc_hd__or2b_1
XFILLER_97_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5108_ _5108_/A _5108_/B vssd1 vssd1 vccd1 vccd1 _5141_/D sky130_fd_sc_hd__nor2_1
XFILLER_85_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6088_ _6088_/A _6185_/A vssd1 vssd1 vccd1 vccd1 _6088_/Y sky130_fd_sc_hd__nor2_1
X_5039_ _5187_/A _5128_/A vssd1 vssd1 vccd1 vccd1 _5211_/B sky130_fd_sc_hd__or2_1
XFILLER_38_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8729_ _8732_/CLK _8729_/D vssd1 vssd1 vccd1 vccd1 _8729_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4410_ _4413_/A vssd1 vssd1 vccd1 vccd1 _4410_/Y sky130_fd_sc_hd__inv_2
X_5390_ _5390_/A vssd1 vssd1 vccd1 vccd1 _8696_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7060_ _7060_/A _7060_/B vssd1 vssd1 vccd1 vccd1 _7061_/B sky130_fd_sc_hd__xor2_1
X_6011_ _6011_/A _6011_/B vssd1 vssd1 vccd1 vccd1 _6027_/A sky130_fd_sc_hd__nor2_1
XFILLER_67_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7962_ _7962_/A _7962_/B vssd1 vssd1 vccd1 vccd1 _7963_/B sky130_fd_sc_hd__and2_1
XFILLER_27_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6913_ _7019_/A _6913_/B vssd1 vssd1 vccd1 vccd1 _7017_/B sky130_fd_sc_hd__xor2_2
X_7893_ _7893_/A vssd1 vssd1 vccd1 vccd1 _7893_/Y sky130_fd_sc_hd__inv_2
XFILLER_62_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6844_ _6846_/A _6846_/B vssd1 vssd1 vccd1 vccd1 _6976_/A sky130_fd_sc_hd__xnor2_1
XFILLER_22_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6775_ _6775_/A _6775_/B vssd1 vssd1 vccd1 vccd1 _6780_/A sky130_fd_sc_hd__xnor2_1
X_8514_ _8514_/A _8514_/B _8514_/C vssd1 vssd1 vccd1 vccd1 _8514_/X sky130_fd_sc_hd__or3_1
X_5726_ _5727_/A _5632_/A _5741_/A vssd1 vssd1 vccd1 vccd1 _5728_/B sky130_fd_sc_hd__a21oi_1
XFILLER_50_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8445_ _8445_/A _8445_/B vssd1 vssd1 vccd1 vccd1 _8471_/A sky130_fd_sc_hd__xnor2_2
X_5657_ _5662_/B _5657_/B vssd1 vssd1 vccd1 vccd1 _5764_/B sky130_fd_sc_hd__xnor2_1
X_8376_ _8376_/A _8378_/C vssd1 vssd1 vccd1 vccd1 _8460_/A sky130_fd_sc_hd__nand2_1
X_5588_ _5688_/A _5725_/B vssd1 vssd1 vccd1 vccd1 _5892_/A sky130_fd_sc_hd__or2_1
X_4608_ _8634_/Q _8633_/Q _8636_/Q _8635_/Q vssd1 vssd1 vccd1 vccd1 _4611_/B sky130_fd_sc_hd__or4_1
X_7327_ _7233_/B _7327_/B vssd1 vssd1 vccd1 vccd1 _7327_/X sky130_fd_sc_hd__and2b_1
X_4539_ _4878_/A vssd1 vssd1 vccd1 vccd1 _4877_/A sky130_fd_sc_hd__clkbuf_1
X_7258_ _7240_/A _7240_/B _7220_/A vssd1 vssd1 vccd1 vccd1 _7350_/A sky130_fd_sc_hd__a21oi_1
XFILLER_89_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6209_ _6209_/A _6209_/B vssd1 vssd1 vccd1 vccd1 _6244_/B sky130_fd_sc_hd__xnor2_1
XFILLER_77_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7189_ _7190_/A _7485_/B vssd1 vssd1 vccd1 vccd1 _7272_/A sky130_fd_sc_hd__and2_1
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4890_ _5272_/B _5156_/A vssd1 vssd1 vccd1 vccd1 _4891_/B sky130_fd_sc_hd__or2_1
XFILLER_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6560_ _6560_/A _6560_/B vssd1 vssd1 vccd1 vccd1 _6560_/Y sky130_fd_sc_hd__nor2_1
X_5511_ _5698_/A _5916_/A vssd1 vssd1 vccd1 vccd1 _5512_/B sky130_fd_sc_hd__nand2_1
XFILLER_8_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6491_ _6491_/A _6491_/B vssd1 vssd1 vccd1 vccd1 _8733_/D sky130_fd_sc_hd__nor2_1
X_8230_ _8228_/Y _8225_/B _8229_/Y vssd1 vssd1 vccd1 vccd1 _8480_/A sky130_fd_sc_hd__a21oi_2
X_5442_ _5440_/C _5436_/Y _5441_/X _5335_/X vssd1 vssd1 vccd1 vccd1 _8706_/D sky130_fd_sc_hd__o211a_1
X_8161_ _8172_/B vssd1 vssd1 vccd1 vccd1 _8514_/B sky130_fd_sc_hd__clkbuf_2
X_5373_ _8691_/Q _5371_/A _5360_/X vssd1 vssd1 vccd1 vccd1 _5374_/B sky130_fd_sc_hd__o21ai_1
X_8092_ _8092_/A _8102_/B vssd1 vssd1 vccd1 vccd1 _8239_/A sky130_fd_sc_hd__nand2_1
X_7112_ _6717_/B _6973_/A _6725_/Y vssd1 vssd1 vccd1 vccd1 _7116_/A sky130_fd_sc_hd__a21o_1
XFILLER_99_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7043_ _7168_/A _7168_/B vssd1 vssd1 vccd1 vccd1 _7165_/B sky130_fd_sc_hd__xor2_1
XFILLER_99_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7945_ _8190_/B vssd1 vssd1 vccd1 vccd1 _8348_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7876_ _8330_/A _8025_/A vssd1 vssd1 vccd1 vccd1 _8103_/A sky130_fd_sc_hd__or2_1
XFILLER_70_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6827_ _7176_/A vssd1 vssd1 vccd1 vccd1 _6966_/B sky130_fd_sc_hd__buf_2
XFILLER_50_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6758_ _6758_/A _6758_/B vssd1 vssd1 vccd1 vccd1 _6758_/Y sky130_fd_sc_hd__nand2_1
X_5709_ _5962_/A _5709_/B vssd1 vssd1 vccd1 vccd1 _5709_/Y sky130_fd_sc_hd__nand2_1
XFILLER_6_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6689_ _7302_/B vssd1 vssd1 vccd1 vccd1 _7050_/A sky130_fd_sc_hd__clkbuf_2
X_8428_ _8428_/A _8428_/B vssd1 vssd1 vccd1 vccd1 _8429_/B sky130_fd_sc_hd__xnor2_1
XFILLER_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8359_ _8353_/X _8487_/B _8358_/Y vssd1 vssd1 vccd1 vccd1 _8360_/B sky130_fd_sc_hd__a21oi_1
XFILLER_104_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_4_12_0_wb_clk_i clkbuf_3_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8783_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_76_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5991_ _5991_/A vssd1 vssd1 vccd1 vccd1 _6183_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7730_ _7821_/A _7752_/B _7729_/X vssd1 vssd1 vccd1 vccd1 _7788_/B sky130_fd_sc_hd__a21o_2
XFILLER_52_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4942_ _4942_/A vssd1 vssd1 vccd1 vccd1 _5153_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_7661_ _7661_/A _7665_/B vssd1 vssd1 vccd1 vccd1 _7662_/B sky130_fd_sc_hd__nand2_1
X_4873_ _4910_/A _4934_/B vssd1 vssd1 vccd1 vccd1 _5033_/A sky130_fd_sc_hd__nor2_1
X_6612_ _8760_/Q _7729_/B vssd1 vssd1 vccd1 vccd1 _6637_/B sky130_fd_sc_hd__xnor2_1
X_7592_ _8780_/Q vssd1 vssd1 vccd1 vccd1 _8593_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6543_ _8765_/Q _6560_/A _6543_/C vssd1 vssd1 vccd1 vccd1 _6543_/X sky130_fd_sc_hd__or3_1
X_6474_ _6478_/C _6474_/B _6517_/B vssd1 vssd1 vccd1 vccd1 _6475_/A sky130_fd_sc_hd__and3b_1
X_8213_ _8496_/S _8239_/A vssd1 vssd1 vccd1 vccd1 _8214_/C sky130_fd_sc_hd__nor2_1
X_5425_ _5617_/A vssd1 vssd1 vccd1 vccd1 _6433_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_99_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8144_ _8135_/A _8135_/B _8143_/X vssd1 vssd1 vccd1 vccd1 _8312_/A sky130_fd_sc_hd__a21o_1
X_5356_ _8685_/Q _8684_/Q _8686_/Q vssd1 vssd1 vccd1 vccd1 _5357_/C sky130_fd_sc_hd__a21o_1
XFILLER_101_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8075_ _7996_/A _8248_/B _8514_/C _7999_/X vssd1 vssd1 vccd1 vccd1 _8181_/B sky130_fd_sc_hd__a31oi_2
X_5287_ _5192_/A _5283_/C _5278_/B _5282_/X _5286_/X vssd1 vssd1 vccd1 vccd1 _5287_/X
+ sky130_fd_sc_hd__o41a_1
XINSDIODE2_5 _5251_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7026_ _6936_/A _6936_/B _6937_/B _7228_/B vssd1 vssd1 vccd1 vccd1 _7223_/A sky130_fd_sc_hd__a22oi_2
XFILLER_95_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8977_ _8977_/A _4472_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[26] sky130_fd_sc_hd__ebufn_8
X_7928_ _7928_/A _7928_/B _7928_/C vssd1 vssd1 vccd1 vccd1 _7929_/B sky130_fd_sc_hd__or3_1
XFILLER_70_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7859_ _7859_/A _7859_/B vssd1 vssd1 vccd1 vccd1 _7860_/B sky130_fd_sc_hd__xnor2_1
XFILLER_51_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5210_ _5210_/A _5210_/B vssd1 vssd1 vccd1 vccd1 _5211_/D sky130_fd_sc_hd__nand2_1
X_6190_ _6190_/A _6190_/B vssd1 vssd1 vccd1 vccd1 _6207_/A sky130_fd_sc_hd__or2_1
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5141_ _5221_/A _5250_/C _5141_/C _5141_/D vssd1 vssd1 vccd1 vccd1 _5141_/X sky130_fd_sc_hd__and4bb_1
XFILLER_69_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5072_ _5096_/B _5069_/X _5071_/X _4818_/A vssd1 vssd1 vccd1 vccd1 _5073_/C sky130_fd_sc_hd__o211a_1
X_8900_ _8900_/A _4381_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[19] sky130_fd_sc_hd__ebufn_8
XFILLER_96_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8762_ _8763_/CLK _8762_/D vssd1 vssd1 vccd1 vccd1 _8762_/Q sky130_fd_sc_hd__dfxtp_1
X_5974_ _5911_/A _5911_/B _5973_/X vssd1 vssd1 vccd1 vccd1 _6055_/A sky130_fd_sc_hd__a21oi_2
X_7713_ _8568_/A _7712_/A _8293_/A _7712_/Y vssd1 vssd1 vccd1 vccd1 _7714_/B sky130_fd_sc_hd__o31a_1
X_4925_ _4925_/A _4925_/B vssd1 vssd1 vccd1 vccd1 _5077_/B sky130_fd_sc_hd__nor2_2
X_8693_ _8704_/CLK _8693_/D vssd1 vssd1 vccd1 vccd1 _8693_/Q sky130_fd_sc_hd__dfxtp_1
X_7644_ _8628_/A vssd1 vssd1 vccd1 vccd1 _7644_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4856_ _5148_/A _4969_/A vssd1 vssd1 vccd1 vccd1 _4856_/Y sky130_fd_sc_hd__nor2_1
XFILLER_20_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7575_ _7575_/A _7575_/B vssd1 vssd1 vccd1 vccd1 _7575_/X sky130_fd_sc_hd__or2_1
X_4787_ _8588_/A _4787_/B vssd1 vssd1 vccd1 vccd1 _4788_/A sky130_fd_sc_hd__and2_1
XFILLER_20_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6526_ _8765_/Q vssd1 vssd1 vccd1 vccd1 _6653_/A sky130_fd_sc_hd__inv_2
XFILLER_4_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6457_ _8728_/Q _6457_/B _8732_/Q _6456_/X vssd1 vssd1 vccd1 vccd1 _7619_/C sky130_fd_sc_hd__or4b_4
X_6388_ _6389_/B _6388_/B vssd1 vssd1 vccd1 vccd1 _6394_/B sky130_fd_sc_hd__and2b_1
X_5408_ _8702_/Q _5408_/B vssd1 vssd1 vccd1 vccd1 _5409_/C sky130_fd_sc_hd__nand2_1
XFILLER_87_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8127_ _8128_/A _8128_/B vssd1 vssd1 vccd1 vccd1 _8222_/A sky130_fd_sc_hd__nand2_2
X_5339_ _8687_/Q _8686_/Q _6535_/A _6532_/B _8689_/Q vssd1 vssd1 vccd1 vccd1 _5339_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_102_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8058_ _8058_/A _8039_/X vssd1 vssd1 vccd1 vccd1 _8145_/B sky130_fd_sc_hd__or2b_1
XFILLER_87_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7009_ _7118_/B _6900_/A _7009_/S vssd1 vssd1 vccd1 vccd1 _7010_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8869__86 vssd1 vssd1 vccd1 vccd1 _8869__86/HI _8978_/A sky130_fd_sc_hd__conb_1
XFILLER_50_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5690_ _6071_/A _5702_/A _5645_/C _6262_/B vssd1 vssd1 vccd1 vccd1 _5704_/B sky130_fd_sc_hd__o211ai_2
XFILLER_61_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4710_ _4946_/A _4732_/B vssd1 vssd1 vccd1 vccd1 _4718_/B sky130_fd_sc_hd__nand2_1
XFILLER_30_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4641_ _8638_/Q _4643_/C _4640_/X vssd1 vssd1 vccd1 vccd1 _4641_/Y sky130_fd_sc_hd__o21ai_1
X_4572_ _6673_/B _4754_/A vssd1 vssd1 vccd1 vccd1 _4702_/A sky130_fd_sc_hd__nand2_1
X_7360_ _7434_/A _7508_/A vssd1 vssd1 vccd1 vccd1 _7360_/Y sky130_fd_sc_hd__nand2_1
X_6311_ _5928_/B _6311_/B _6311_/C vssd1 vssd1 vccd1 vccd1 _6313_/A sky130_fd_sc_hd__and3b_1
X_7291_ _7291_/A _7291_/B vssd1 vssd1 vccd1 vccd1 _7292_/B sky130_fd_sc_hd__nand2_1
X_6242_ _6242_/A _6342_/A vssd1 vssd1 vccd1 vccd1 _6286_/A sky130_fd_sc_hd__xnor2_1
XFILLER_89_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6173_ _6173_/A _6230_/B vssd1 vssd1 vccd1 vccd1 _6302_/B sky130_fd_sc_hd__xor2_2
XFILLER_69_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5124_ _5275_/B _5184_/B _5148_/B _5124_/D vssd1 vssd1 vccd1 vccd1 _5124_/X sky130_fd_sc_hd__or4_1
X_5055_ _5277_/B _5225_/B _5228_/A _5055_/D vssd1 vssd1 vccd1 vccd1 _5055_/X sky130_fd_sc_hd__or4_1
XFILLER_84_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5957_ _5957_/A _5957_/B vssd1 vssd1 vccd1 vccd1 _6128_/B sky130_fd_sc_hd__xor2_2
X_8745_ _8765_/CLK _8745_/D vssd1 vssd1 vccd1 vccd1 _8745_/Q sky130_fd_sc_hd__dfxtp_1
X_8676_ _8776_/CLK _8676_/D vssd1 vssd1 vccd1 vccd1 _8676_/Q sky130_fd_sc_hd__dfxtp_1
X_4908_ _4910_/A vssd1 vssd1 vccd1 vccd1 _5040_/B sky130_fd_sc_hd__clkbuf_2
X_5888_ _5888_/A _5888_/B vssd1 vssd1 vccd1 vccd1 _5973_/B sky130_fd_sc_hd__nand2_1
X_7627_ _7649_/B vssd1 vssd1 vccd1 vccd1 _7627_/X sky130_fd_sc_hd__buf_2
XFILLER_21_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4839_ _4916_/B vssd1 vssd1 vccd1 vccd1 _5032_/B sky130_fd_sc_hd__inv_2
X_7558_ _7558_/A _7558_/B vssd1 vssd1 vccd1 vccd1 _7559_/B sky130_fd_sc_hd__nand2_1
X_7489_ _7489_/A _7489_/B vssd1 vssd1 vccd1 vccd1 _7489_/Y sky130_fd_sc_hd__nor2_1
X_6509_ _6509_/A vssd1 vssd1 vccd1 vccd1 _8739_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6860_ _7489_/A _6834_/B _6858_/C vssd1 vssd1 vccd1 vccd1 _6861_/B sky130_fd_sc_hd__a21oi_1
XFILLER_19_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5811_ _5811_/A _5811_/B _5811_/C vssd1 vssd1 vccd1 vccd1 _5811_/X sky130_fd_sc_hd__and3_1
X_6791_ _6835_/A vssd1 vssd1 vccd1 vccd1 _6792_/B sky130_fd_sc_hd__clkbuf_2
X_8530_ _7913_/A _7917_/A _8382_/B _7800_/Y vssd1 vssd1 vccd1 vccd1 _8531_/B sky130_fd_sc_hd__o211a_1
X_5742_ _6081_/A _5827_/A _5741_/Y vssd1 vssd1 vccd1 vccd1 _5743_/B sky130_fd_sc_hd__a21oi_1
XFILLER_34_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8461_ _7999_/X _8460_/Y _8461_/S vssd1 vssd1 vccd1 vccd1 _8513_/B sky130_fd_sc_hd__mux2_1
X_5673_ _5673_/A _5673_/B vssd1 vssd1 vccd1 vccd1 _5674_/C sky130_fd_sc_hd__and2_1
X_8392_ _8277_/A _8277_/B _8272_/C vssd1 vssd1 vccd1 vccd1 _8457_/B sky130_fd_sc_hd__a21o_1
X_7412_ _7412_/A _7412_/B vssd1 vssd1 vccd1 vccd1 _7415_/A sky130_fd_sc_hd__xnor2_1
X_4624_ _4631_/C _4679_/A _4624_/C vssd1 vssd1 vccd1 vccd1 _4625_/A sky130_fd_sc_hd__and3b_1
X_7343_ _7350_/A _7350_/B vssd1 vssd1 vccd1 vccd1 _7344_/B sky130_fd_sc_hd__xor2_1
X_4555_ _5231_/A vssd1 vssd1 vccd1 vccd1 _4555_/X sky130_fd_sc_hd__clkbuf_2
X_7274_ _7274_/A vssd1 vssd1 vccd1 vccd1 _7501_/A sky130_fd_sc_hd__clkbuf_2
X_4486_ _4486_/A vssd1 vssd1 vccd1 vccd1 _4486_/Y sky130_fd_sc_hd__inv_2
X_6225_ _6152_/A _6152_/B _6224_/X vssd1 vssd1 vccd1 vccd1 _6234_/A sky130_fd_sc_hd__a21o_1
X_6156_ _6156_/A _6156_/B vssd1 vssd1 vccd1 vccd1 _6158_/A sky130_fd_sc_hd__nand2_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5107_ _5107_/A _5107_/B vssd1 vssd1 vccd1 vccd1 _5117_/B sky130_fd_sc_hd__nand2_2
X_6087_ _6087_/A _6087_/B vssd1 vssd1 vccd1 vccd1 _6099_/A sky130_fd_sc_hd__xnor2_2
XFILLER_57_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5038_ _5038_/A _5038_/B vssd1 vssd1 vccd1 vccd1 _5038_/X sky130_fd_sc_hd__or2_1
XFILLER_65_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6989_ _7069_/A _7069_/B vssd1 vssd1 vccd1 vccd1 _7067_/C sky130_fd_sc_hd__nand2_1
XFILLER_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8728_ _8730_/CLK _8728_/D vssd1 vssd1 vccd1 vccd1 _8728_/Q sky130_fd_sc_hd__dfxtp_1
X_8659_ _8778_/CLK _8659_/D vssd1 vssd1 vccd1 vccd1 _8659_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8839__56 vssd1 vssd1 vccd1 vccd1 _8839__56/HI _8948_/A sky130_fd_sc_hd__conb_1
XFILLER_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6010_ _6055_/A _6055_/B vssd1 vssd1 vccd1 vccd1 _6029_/A sky130_fd_sc_hd__xor2_1
XFILLER_98_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8853__70 vssd1 vssd1 vccd1 vccd1 _8853__70/HI _8962_/A sky130_fd_sc_hd__conb_1
XFILLER_79_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7961_ _7962_/A _7962_/B vssd1 vssd1 vccd1 vccd1 _8056_/A sky130_fd_sc_hd__nor2_1
XFILLER_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7892_ _7892_/A _7892_/B vssd1 vssd1 vccd1 vccd1 _7892_/X sky130_fd_sc_hd__or2_1
X_6912_ _6910_/X _6912_/B vssd1 vssd1 vccd1 vccd1 _6913_/B sky130_fd_sc_hd__and2b_1
XFILLER_62_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6843_ _6848_/A _6848_/B vssd1 vssd1 vccd1 vccd1 _6846_/B sky130_fd_sc_hd__xnor2_1
XFILLER_35_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6774_ _6774_/A vssd1 vssd1 vccd1 vccd1 _7118_/B sky130_fd_sc_hd__buf_2
X_8513_ _8513_/A _8513_/B vssd1 vssd1 vccd1 vccd1 _8513_/Y sky130_fd_sc_hd__nand2_1
X_5725_ _5725_/A _5725_/B vssd1 vssd1 vccd1 vccd1 _5741_/A sky130_fd_sc_hd__nor2_1
XFILLER_50_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8444_ _8442_/X _8444_/B vssd1 vssd1 vccd1 vccd1 _8445_/B sky130_fd_sc_hd__and2b_1
X_5656_ _5666_/A _5766_/C vssd1 vssd1 vccd1 vccd1 _5657_/B sky130_fd_sc_hd__xnor2_1
X_4607_ _8632_/Q _8631_/Q vssd1 vssd1 vccd1 vccd1 _4620_/A sky130_fd_sc_hd__or2_1
X_8375_ _8280_/A _8280_/B _8280_/D _8374_/Y vssd1 vssd1 vccd1 vccd1 _8396_/A sky130_fd_sc_hd__a31o_1
X_5587_ _5587_/A _5587_/B vssd1 vssd1 vccd1 vccd1 _5725_/B sky130_fd_sc_hd__xnor2_1
XFILLER_104_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7326_ _7216_/A _7216_/B _7325_/X vssd1 vssd1 vccd1 vccd1 _7340_/A sky130_fd_sc_hd__a21o_1
X_4538_ _7672_/B vssd1 vssd1 vccd1 vccd1 _4878_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_89_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4469_ _4481_/A vssd1 vssd1 vccd1 vccd1 _4474_/A sky130_fd_sc_hd__clkbuf_2
X_7257_ _7257_/A _7257_/B vssd1 vssd1 vccd1 vccd1 _7344_/A sky130_fd_sc_hd__nand2_1
X_6208_ _6208_/A _6208_/B vssd1 vssd1 vccd1 vccd1 _6209_/B sky130_fd_sc_hd__nor2_1
X_7188_ _7204_/A vssd1 vssd1 vccd1 vccd1 _7485_/B sky130_fd_sc_hd__buf_2
X_6139_ _6064_/A _6064_/B _6065_/B _6065_/A vssd1 vssd1 vccd1 vccd1 _6161_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_58_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5510_ _5530_/A _5530_/B vssd1 vssd1 vccd1 vccd1 _5916_/A sky130_fd_sc_hd__xnor2_4
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6490_ _8733_/Q _6492_/C _6483_/X vssd1 vssd1 vccd1 vccd1 _6491_/B sky130_fd_sc_hd__o21ai_1
X_5441_ _5477_/B _5440_/X vssd1 vssd1 vccd1 vccd1 _5441_/X sky130_fd_sc_hd__or2b_1
X_8160_ _8272_/A _8272_/B vssd1 vssd1 vccd1 vccd1 _8169_/A sky130_fd_sc_hd__or2_1
X_5372_ _8691_/Q _8690_/Q _5372_/C vssd1 vssd1 vccd1 vccd1 _5377_/C sky130_fd_sc_hd__and3_1
X_8091_ _8355_/A vssd1 vssd1 vccd1 vccd1 _8336_/A sky130_fd_sc_hd__clkbuf_2
X_7111_ _7111_/A _7111_/B vssd1 vssd1 vccd1 vccd1 _7116_/B sky130_fd_sc_hd__xnor2_1
XFILLER_86_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7042_ _7223_/A _7042_/B vssd1 vssd1 vccd1 vccd1 _7168_/B sky130_fd_sc_hd__xnor2_1
XFILLER_82_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7944_ _7843_/B _7845_/B _7943_/Y vssd1 vssd1 vccd1 vccd1 _8190_/B sky130_fd_sc_hd__a21o_1
XFILLER_55_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7875_ _7875_/A _7875_/B vssd1 vssd1 vccd1 vccd1 _7888_/A sky130_fd_sc_hd__nor2_1
XFILLER_23_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6826_ _7020_/B vssd1 vssd1 vccd1 vccd1 _7176_/A sky130_fd_sc_hd__buf_2
XFILLER_50_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6757_ _6757_/A _6757_/B _6757_/C vssd1 vssd1 vccd1 vccd1 _6866_/D sky130_fd_sc_hd__or3_1
X_5708_ _6398_/A _5711_/A vssd1 vssd1 vccd1 vccd1 _5709_/B sky130_fd_sc_hd__nand2_1
XFILLER_6_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6688_ _6688_/A vssd1 vssd1 vccd1 vccd1 _7302_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_8427_ _8427_/A _8427_/B vssd1 vssd1 vccd1 vccd1 _8428_/B sky130_fd_sc_hd__xor2_1
X_5639_ _6378_/C _6197_/A _5639_/C vssd1 vssd1 vccd1 vccd1 _5640_/B sky130_fd_sc_hd__nor3_1
X_8358_ _8358_/A _8358_/B vssd1 vssd1 vccd1 vccd1 _8358_/Y sky130_fd_sc_hd__nor2_1
XFILLER_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8809__26 vssd1 vssd1 vccd1 vccd1 _8809__26/HI _8904_/A sky130_fd_sc_hd__conb_1
X_7309_ _7309_/A _7309_/B vssd1 vssd1 vccd1 vccd1 _7390_/A sky130_fd_sc_hd__nand2_1
X_8289_ _8568_/B _8289_/B vssd1 vssd1 vccd1 vccd1 _8505_/A sky130_fd_sc_hd__nand2_1
XFILLER_104_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8823__40 vssd1 vssd1 vccd1 vccd1 _8823__40/HI _8918_/A sky130_fd_sc_hd__conb_1
XFILLER_83_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5990_ _6068_/A _6068_/B vssd1 vssd1 vccd1 vccd1 _5996_/A sky130_fd_sc_hd__nand2_1
X_4941_ _5209_/A _5272_/C vssd1 vssd1 vccd1 vccd1 _4957_/A sky130_fd_sc_hd__or2_1
XFILLER_45_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7660_ _7775_/A _8767_/Q vssd1 vssd1 vccd1 vccd1 _7665_/B sky130_fd_sc_hd__or2_1
X_4872_ _4878_/B _4872_/B _4762_/A _4877_/A vssd1 vssd1 vccd1 vccd1 _4934_/B sky130_fd_sc_hd__or4bb_2
X_6611_ _6648_/A _6648_/B vssd1 vssd1 vccd1 vccd1 _7309_/A sky130_fd_sc_hd__nand2_4
X_7591_ _8781_/Q vssd1 vssd1 vccd1 vccd1 _7734_/A sky130_fd_sc_hd__clkbuf_2
X_6542_ _7562_/A _7556_/A _8762_/Q vssd1 vssd1 vccd1 vccd1 _6543_/C sky130_fd_sc_hd__o21a_1
XFILLER_9_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6473_ _8728_/Q _6473_/B vssd1 vssd1 vccd1 vccd1 _6474_/B sky130_fd_sc_hd__or2_1
X_8212_ _8358_/A vssd1 vssd1 vccd1 vccd1 _8496_/S sky130_fd_sc_hd__clkbuf_2
X_5424_ _8724_/Q vssd1 vssd1 vccd1 vccd1 _5617_/A sky130_fd_sc_hd__inv_2
X_8143_ _8134_/B _8143_/B vssd1 vssd1 vccd1 vccd1 _8143_/X sky130_fd_sc_hd__and2b_1
X_5355_ _5355_/A vssd1 vssd1 vccd1 vccd1 _5389_/B sky130_fd_sc_hd__buf_2
XFILLER_101_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8074_ _8261_/A _8376_/A vssd1 vssd1 vccd1 vccd1 _8514_/C sky130_fd_sc_hd__nand2_1
X_5286_ _5286_/A _5286_/B vssd1 vssd1 vccd1 vccd1 _5286_/X sky130_fd_sc_hd__or2_1
XINSDIODE2_6 _5226_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7025_ _7025_/A _7167_/A vssd1 vssd1 vccd1 vccd1 _7168_/A sky130_fd_sc_hd__xnor2_1
XFILLER_28_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8976_ _8976_/A _4471_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[25] sky130_fd_sc_hd__ebufn_8
XFILLER_82_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7927_ _7928_/A _7928_/B _7928_/C vssd1 vssd1 vccd1 vccd1 _8018_/A sky130_fd_sc_hd__o21a_1
XFILLER_70_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7858_ _7858_/A _7858_/B vssd1 vssd1 vccd1 vccd1 _7859_/B sky130_fd_sc_hd__nor2_1
X_6809_ _6809_/A _6897_/A vssd1 vssd1 vccd1 vccd1 _6856_/A sky130_fd_sc_hd__or2_1
XFILLER_23_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7789_ _7789_/A _7789_/B vssd1 vssd1 vccd1 vccd1 _7899_/A sky130_fd_sc_hd__xor2_1
XFILLER_11_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5140_ _5197_/D vssd1 vssd1 vccd1 vccd1 _5140_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5071_ _5168_/A _5201_/B _5071_/C _5071_/D vssd1 vssd1 vccd1 vccd1 _5071_/X sky130_fd_sc_hd__or4_1
XFILLER_49_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5973_ _5906_/B _5973_/B vssd1 vssd1 vccd1 vccd1 _5973_/X sky130_fd_sc_hd__and2b_1
XFILLER_64_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8761_ _8763_/CLK _8761_/D vssd1 vssd1 vccd1 vccd1 _8761_/Q sky130_fd_sc_hd__dfxtp_1
X_7712_ _7712_/A _7764_/A vssd1 vssd1 vccd1 vccd1 _7712_/Y sky130_fd_sc_hd__nand2_1
XFILLER_52_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4924_ _5206_/A _4978_/A vssd1 vssd1 vccd1 vccd1 _5062_/A sky130_fd_sc_hd__or2_1
X_8692_ _8704_/CLK _8692_/D vssd1 vssd1 vccd1 vccd1 _8692_/Q sky130_fd_sc_hd__dfxtp_1
X_7643_ _7637_/A _7627_/X _7641_/X _7642_/X vssd1 vssd1 vccd1 vccd1 _8770_/D sky130_fd_sc_hd__o211a_1
XFILLER_20_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4855_ _5206_/B vssd1 vssd1 vccd1 vccd1 _4969_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_33_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7574_ _7575_/A _7575_/B vssd1 vssd1 vccd1 vccd1 _7586_/S sky130_fd_sc_hd__nand2_1
X_4786_ _4767_/B _5040_/A _4785_/X _5315_/A _4541_/X vssd1 vssd1 vccd1 vccd1 _4787_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_20_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6525_ _6525_/A vssd1 vssd1 vccd1 vccd1 _8745_/D sky130_fd_sc_hd__clkbuf_1
X_6456_ _8744_/Q _6456_/B _8745_/Q _8743_/Q vssd1 vssd1 vccd1 vccd1 _6456_/X sky130_fd_sc_hd__and4b_1
X_6387_ _7656_/B vssd1 vssd1 vccd1 vccd1 _6387_/X sky130_fd_sc_hd__clkbuf_2
X_5407_ _8702_/Q _5408_/B vssd1 vssd1 vccd1 vccd1 _5409_/B sky130_fd_sc_hd__or2_1
X_8126_ _8304_/A _8126_/B vssd1 vssd1 vccd1 vccd1 _8128_/B sky130_fd_sc_hd__nor2_1
X_5338_ _8688_/Q vssd1 vssd1 vccd1 vccd1 _6532_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_102_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8057_ _8057_/A _8057_/B vssd1 vssd1 vccd1 vccd1 _8143_/B sky130_fd_sc_hd__nand2_1
X_7008_ _6760_/X _6758_/Y _6759_/X _6784_/B _6752_/A vssd1 vssd1 vccd1 vccd1 _7009_/S
+ sky130_fd_sc_hd__a311o_1
X_5269_ _5269_/A _5285_/B vssd1 vssd1 vccd1 vccd1 _5291_/B sky130_fd_sc_hd__or2_1
XFILLER_47_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8959_ _8959_/A _4446_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[8] sky130_fd_sc_hd__ebufn_8
XFILLER_43_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4640_ _4640_/A vssd1 vssd1 vccd1 vccd1 _4640_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_30_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6310_ _6232_/A _6232_/B _6309_/X vssd1 vssd1 vccd1 vccd1 _6314_/A sky130_fd_sc_hd__a21o_1
X_4571_ _4814_/A _4814_/B _4571_/C _4692_/C vssd1 vssd1 vccd1 vccd1 _4573_/B sky130_fd_sc_hd__or4_1
X_7290_ _7291_/A _7291_/B vssd1 vssd1 vccd1 vccd1 _7290_/Y sky130_fd_sc_hd__nor2_1
X_6241_ _6107_/B _6160_/B _6240_/Y vssd1 vssd1 vccd1 vccd1 _6342_/A sky130_fd_sc_hd__a21oi_2
X_6172_ _6172_/A _6252_/B vssd1 vssd1 vccd1 vccd1 _6230_/B sky130_fd_sc_hd__and2_1
X_5123_ _5123_/A _5187_/A _5184_/B vssd1 vssd1 vccd1 vccd1 _5123_/X sky130_fd_sc_hd__or3_1
XFILLER_69_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5054_ _5135_/A _5054_/B _5054_/C _5124_/D vssd1 vssd1 vccd1 vccd1 _5055_/D sky130_fd_sc_hd__or4_1
XFILLER_38_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5956_ _5967_/B _5956_/B vssd1 vssd1 vccd1 vccd1 _5957_/B sky130_fd_sc_hd__xnor2_1
XFILLER_40_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8744_ _8765_/CLK _8744_/D vssd1 vssd1 vccd1 vccd1 _8744_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5887_ _5887_/A _5887_/B vssd1 vssd1 vccd1 vccd1 _5971_/A sky130_fd_sc_hd__nand2_1
X_8675_ _8776_/CLK _8675_/D vssd1 vssd1 vccd1 vccd1 _8675_/Q sky130_fd_sc_hd__dfxtp_1
X_4907_ _5154_/A _5179_/B vssd1 vssd1 vccd1 vccd1 _4920_/A sky130_fd_sc_hd__or2_1
XFILLER_40_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7626_ _8768_/Q _8609_/A _7625_/Y vssd1 vssd1 vccd1 vccd1 _8768_/D sky130_fd_sc_hd__a21oi_1
X_4838_ _4774_/A _4878_/C _4878_/A _4878_/B vssd1 vssd1 vccd1 vccd1 _4916_/B sky130_fd_sc_hd__and4b_1
X_7557_ _7558_/A _7558_/B vssd1 vssd1 vccd1 vccd1 _7557_/Y sky130_fd_sc_hd__nor2_1
X_4769_ _4769_/A vssd1 vssd1 vccd1 vccd1 _8662_/D sky130_fd_sc_hd__clkbuf_1
X_7488_ _7423_/A _7423_/B _7487_/Y vssd1 vssd1 vccd1 vccd1 _7500_/A sky130_fd_sc_hd__a21o_1
X_6508_ _6510_/B _6508_/B _6508_/C vssd1 vssd1 vccd1 vccd1 _6509_/A sky130_fd_sc_hd__and3b_1
X_6439_ _8740_/Q _8742_/Q _8741_/Q _8739_/Q vssd1 vssd1 vccd1 vccd1 _6456_/B sky130_fd_sc_hd__and4bb_1
XFILLER_0_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8109_ _8109_/A _8236_/C vssd1 vssd1 vccd1 vccd1 _8487_/A sky130_fd_sc_hd__xnor2_4
XFILLER_102_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5810_ _5810_/A _5810_/B _5810_/C vssd1 vssd1 vccd1 vccd1 _5810_/X sky130_fd_sc_hd__and3_1
X_6790_ _6866_/D vssd1 vssd1 vccd1 vccd1 _6836_/A sky130_fd_sc_hd__clkbuf_2
X_5741_ _5741_/A _5751_/A vssd1 vssd1 vccd1 vccd1 _5741_/Y sky130_fd_sc_hd__nor2_1
XFILLER_22_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8460_ _8460_/A vssd1 vssd1 vccd1 vccd1 _8460_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5672_ _5673_/A _5673_/B vssd1 vssd1 vccd1 vccd1 _5715_/A sky130_fd_sc_hd__nor2_1
X_7411_ _7411_/A _7411_/B vssd1 vssd1 vccd1 vccd1 _7412_/B sky130_fd_sc_hd__nor2_1
XFILLER_30_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8391_ _8463_/B _8463_/C vssd1 vssd1 vccd1 vccd1 _8393_/A sky130_fd_sc_hd__xnor2_2
X_4623_ _8632_/Q _8631_/Q _8633_/Q vssd1 vssd1 vccd1 vccd1 _4624_/C sky130_fd_sc_hd__a21o_1
X_7342_ _7342_/A _7342_/B vssd1 vssd1 vccd1 vccd1 _7350_/B sky130_fd_sc_hd__xnor2_2
X_4554_ _4733_/B vssd1 vssd1 vccd1 vccd1 _5231_/A sky130_fd_sc_hd__clkbuf_2
X_7273_ _7409_/B _7272_/C _7272_/A vssd1 vssd1 vccd1 vccd1 _7276_/B sky130_fd_sc_hd__a21o_1
XFILLER_103_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4485_ _4486_/A vssd1 vssd1 vccd1 vccd1 _4485_/Y sky130_fd_sc_hd__inv_2
X_6224_ _6224_/A _6224_/B vssd1 vssd1 vccd1 vccd1 _6224_/X sky130_fd_sc_hd__and2_1
XFILLER_103_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6155_ _6155_/A _6235_/A vssd1 vssd1 vccd1 vccd1 _6159_/A sky130_fd_sc_hd__xor2_1
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6086_ _6181_/A _6181_/B vssd1 vssd1 vccd1 vccd1 _6087_/B sky130_fd_sc_hd__xnor2_2
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5106_ _8654_/Q vssd1 vssd1 vccd1 vccd1 _5160_/A sky130_fd_sc_hd__inv_2
X_5037_ _5188_/A _5285_/A _5159_/D _5215_/C vssd1 vssd1 vccd1 vccd1 _5038_/B sky130_fd_sc_hd__or4_1
XFILLER_53_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6988_ _6988_/A _6988_/B vssd1 vssd1 vccd1 vccd1 _7069_/B sky130_fd_sc_hd__xnor2_1
X_8727_ _8765_/CLK _8727_/D vssd1 vssd1 vccd1 vccd1 _8727_/Q sky130_fd_sc_hd__dfxtp_1
X_5939_ _5939_/A _5939_/B vssd1 vssd1 vccd1 vccd1 _5940_/B sky130_fd_sc_hd__xnor2_1
XFILLER_40_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8658_ _8778_/CLK _8658_/D vssd1 vssd1 vccd1 vccd1 _8658_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_21_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7609_ _8767_/Q vssd1 vssd1 vccd1 vccd1 _7637_/B sky130_fd_sc_hd__inv_2
X_8589_ _7624_/X _8573_/X _8587_/X _8588_/Y vssd1 vssd1 vccd1 vccd1 _8778_/D sky130_fd_sc_hd__a31oi_1
XFILLER_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7960_ _7860_/A _7860_/B _7959_/Y vssd1 vssd1 vccd1 vccd1 _7962_/B sky130_fd_sc_hd__a21oi_1
XFILLER_67_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7891_ _7891_/A _7891_/B vssd1 vssd1 vccd1 vccd1 _7976_/B sky130_fd_sc_hd__or2_1
X_6911_ _6866_/D _6910_/A _6910_/B _6910_/C vssd1 vssd1 vccd1 vccd1 _6912_/B sky130_fd_sc_hd__a31o_1
X_6842_ _6881_/A _6881_/B vssd1 vssd1 vccd1 vccd1 _6848_/B sky130_fd_sc_hd__xor2_1
XFILLER_50_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6773_ _6775_/A _6775_/B vssd1 vssd1 vccd1 vccd1 _7400_/B sky130_fd_sc_hd__xor2_4
X_8512_ _8512_/A _8512_/B vssd1 vssd1 vccd1 vccd1 _8536_/A sky130_fd_sc_hd__nor2_1
X_5724_ _5891_/A _5819_/C _5819_/D vssd1 vssd1 vccd1 vccd1 _5835_/A sky130_fd_sc_hd__or3_2
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8443_ _8443_/A _8443_/B _8441_/Y vssd1 vssd1 vccd1 vccd1 _8444_/B sky130_fd_sc_hd__or3b_1
X_5655_ _5853_/A _5655_/B vssd1 vssd1 vccd1 vccd1 _5766_/C sky130_fd_sc_hd__nor2_2
X_8374_ _8279_/A _8279_/B _8279_/C vssd1 vssd1 vccd1 vccd1 _8374_/Y sky130_fd_sc_hd__a21oi_1
X_4606_ _8638_/Q _8637_/Q _8640_/Q _4606_/D vssd1 vssd1 vccd1 vccd1 _4612_/B sky130_fd_sc_hd__or4_1
X_5586_ _5585_/A _5585_/B _5564_/A vssd1 vssd1 vccd1 vccd1 _5587_/A sky130_fd_sc_hd__a21o_1
X_7325_ _7215_/B _7325_/B vssd1 vssd1 vccd1 vccd1 _7325_/X sky130_fd_sc_hd__and2b_1
XFILLER_89_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4537_ _6621_/B vssd1 vssd1 vccd1 vccd1 _7672_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_104_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4468_ _4468_/A vssd1 vssd1 vccd1 vccd1 _4468_/Y sky130_fd_sc_hd__inv_2
X_7256_ _7256_/A _7239_/B vssd1 vssd1 vccd1 vccd1 _7257_/B sky130_fd_sc_hd__or2b_1
XFILLER_89_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6207_ _6207_/A _6207_/B _6207_/C vssd1 vssd1 vccd1 vccd1 _6208_/B sky130_fd_sc_hd__and3_1
XFILLER_77_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7187_ _7011_/A _6912_/B _7186_/X _6910_/X vssd1 vssd1 vccd1 vccd1 _7204_/A sky130_fd_sc_hd__a211o_1
X_6138_ _6123_/A _6123_/B _6137_/Y vssd1 vssd1 vccd1 vccd1 _6217_/B sky130_fd_sc_hd__a21o_1
XFILLER_100_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4399_ _4400_/A vssd1 vssd1 vccd1 vccd1 _4399_/Y sky130_fd_sc_hd__inv_2
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6069_ _6192_/B vssd1 vssd1 vccd1 vccd1 _6264_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_81_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5440_ _5478_/A _5484_/A _5440_/C _5440_/D vssd1 vssd1 vccd1 vccd1 _5440_/X sky130_fd_sc_hd__or4_1
XFILLER_8_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5371_ _5371_/A _5371_/B vssd1 vssd1 vccd1 vccd1 _8690_/D sky130_fd_sc_hd__nor2_1
X_8090_ _8330_/B vssd1 vssd1 vccd1 vccd1 _8355_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7110_ _7110_/A _7110_/B vssd1 vssd1 vccd1 vccd1 _7111_/B sky130_fd_sc_hd__xnor2_1
X_7041_ _7041_/A _7041_/B vssd1 vssd1 vccd1 vccd1 _7042_/B sky130_fd_sc_hd__xor2_1
XFILLER_67_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7943_ _7943_/A _7943_/B vssd1 vssd1 vccd1 vccd1 _7943_/Y sky130_fd_sc_hd__nor2_1
XFILLER_67_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7874_ _7872_/B _7773_/C _7773_/A vssd1 vssd1 vccd1 vccd1 _7875_/B sky130_fd_sc_hd__o21a_1
Xclkbuf_3_7_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
X_6825_ _6825_/A _7416_/A vssd1 vssd1 vccd1 vccd1 _6973_/A sky130_fd_sc_hd__nor2_2
X_6756_ _6775_/A _6775_/B _6755_/X vssd1 vssd1 vccd1 vccd1 _6757_/C sky130_fd_sc_hd__a21oi_2
X_5707_ _6398_/A _5711_/A vssd1 vssd1 vccd1 vccd1 _5962_/A sky130_fd_sc_hd__or2_1
X_6687_ _7030_/A vssd1 vssd1 vccd1 vccd1 _6809_/A sky130_fd_sc_hd__clkbuf_2
X_8426_ _8337_/A _8337_/B _8425_/X vssd1 vssd1 vccd1 vccd1 _8427_/B sky130_fd_sc_hd__a21oi_1
X_5638_ _6068_/B _6193_/A vssd1 vssd1 vccd1 vccd1 _5639_/C sky130_fd_sc_hd__nor2_1
X_8357_ _8357_/A _8420_/B vssd1 vssd1 vccd1 vccd1 _8487_/B sky130_fd_sc_hd__xnor2_2
X_5569_ _5680_/A _5680_/B _5568_/X vssd1 vssd1 vccd1 vccd1 _5585_/B sky130_fd_sc_hd__a21o_2
XFILLER_88_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7308_ _7397_/A _7397_/B vssd1 vssd1 vccd1 vccd1 _7316_/A sky130_fd_sc_hd__xor2_1
XFILLER_2_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8288_ _8428_/A _8288_/B vssd1 vssd1 vccd1 vccd1 _8340_/A sky130_fd_sc_hd__nand2_1
X_7239_ _7256_/A _7239_/B vssd1 vssd1 vccd1 vccd1 _7240_/B sky130_fd_sc_hd__xnor2_1
XFILLER_77_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4940_ _4956_/A _5201_/A _5201_/B vssd1 vssd1 vccd1 vccd1 _5272_/C sky130_fd_sc_hd__nor3_4
X_4871_ _4892_/A vssd1 vssd1 vccd1 vccd1 _4910_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7590_ _7590_/A vssd1 vssd1 vccd1 vccd1 _8765_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6610_ _7558_/A _7739_/B vssd1 vssd1 vccd1 vccd1 _6648_/B sky130_fd_sc_hd__nand2_1
X_6541_ _7562_/A _7556_/A _8759_/Q _7578_/B _8762_/Q vssd1 vssd1 vccd1 vccd1 _6541_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_9_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6472_ _8728_/Q _6473_/B vssd1 vssd1 vccd1 vccd1 _6478_/C sky130_fd_sc_hd__and2_1
X_8211_ _8428_/A _8288_/B vssd1 vssd1 vccd1 vccd1 _8214_/B sky130_fd_sc_hd__xor2_1
X_5423_ _8724_/Q _5440_/C _5417_/X _5422_/X vssd1 vssd1 vccd1 vccd1 _5423_/X sky130_fd_sc_hd__o31a_1
X_8142_ _8556_/A _8559_/B _8556_/B vssd1 vssd1 vccd1 vccd1 _8562_/C sky130_fd_sc_hd__a21bo_1
X_5354_ _8686_/Q _8685_/Q _8684_/Q vssd1 vssd1 vccd1 vccd1 _5359_/B sky130_fd_sc_hd__and3_1
XFILLER_87_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8073_ _8073_/A vssd1 vssd1 vccd1 vccd1 _8248_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_59_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5285_ _5285_/A _5285_/B _5285_/C _5285_/D vssd1 vssd1 vccd1 vccd1 _5286_/B sky130_fd_sc_hd__or4_1
XINSDIODE2_7 _5240_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7024_ _7024_/A _7024_/B vssd1 vssd1 vccd1 vccd1 _7167_/A sky130_fd_sc_hd__xnor2_1
XFILLER_28_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8975_ _8975_/A _4470_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[24] sky130_fd_sc_hd__ebufn_8
X_7926_ _8008_/A _8376_/A vssd1 vssd1 vccd1 vccd1 _7928_/C sky130_fd_sc_hd__xnor2_1
XFILLER_82_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7857_ _7856_/B _7938_/A vssd1 vssd1 vccd1 vccd1 _7858_/B sky130_fd_sc_hd__and2b_1
XFILLER_23_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6808_ _6963_/A _6845_/B _6807_/X vssd1 vssd1 vccd1 vccd1 _6823_/A sky130_fd_sc_hd__a21o_1
X_7788_ _7788_/A _7788_/B vssd1 vssd1 vccd1 vccd1 _7904_/A sky130_fd_sc_hd__xor2_4
XFILLER_23_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6739_ _8752_/Q _7700_/A vssd1 vssd1 vccd1 vccd1 _6755_/B sky130_fd_sc_hd__and2b_2
XFILLER_23_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8409_ _8344_/A _8409_/B vssd1 vssd1 vccd1 vccd1 _8409_/X sky130_fd_sc_hd__and2b_1
XFILLER_74_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5070_ _5274_/B _5036_/B _5145_/B vssd1 vssd1 vccd1 vccd1 _5071_/D sky130_fd_sc_hd__o21a_1
XFILLER_84_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5972_ _5940_/A _5940_/B _5971_/Y vssd1 vssd1 vccd1 vccd1 _6053_/A sky130_fd_sc_hd__a21boi_1
XFILLER_92_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8760_ _8763_/CLK _8760_/D vssd1 vssd1 vccd1 vccd1 _8760_/Q sky130_fd_sc_hd__dfxtp_1
X_7711_ _7711_/A _7710_/X vssd1 vssd1 vccd1 vccd1 _7764_/A sky130_fd_sc_hd__or2b_1
XFILLER_18_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4923_ _5148_/B _5077_/C vssd1 vssd1 vccd1 vccd1 _4978_/A sky130_fd_sc_hd__or2_1
X_8691_ _8704_/CLK _8691_/D vssd1 vssd1 vccd1 vccd1 _8691_/Q sky130_fd_sc_hd__dfxtp_1
X_4854_ _5159_/D _5050_/D vssd1 vssd1 vccd1 vccd1 _5206_/B sky130_fd_sc_hd__or2_1
X_7642_ _7642_/A vssd1 vssd1 vccd1 vccd1 _7642_/X sky130_fd_sc_hd__clkbuf_2
X_4785_ _4549_/A _4897_/B _5100_/A _4541_/X vssd1 vssd1 vccd1 vccd1 _4785_/X sky130_fd_sc_hd__a31o_1
X_7573_ _6660_/A _7579_/B _7572_/X vssd1 vssd1 vccd1 vccd1 _7575_/B sky130_fd_sc_hd__a21oi_1
X_6524_ _6522_/Y _6524_/B vssd1 vssd1 vccd1 vccd1 _6525_/A sky130_fd_sc_hd__and2b_1
X_6455_ _8726_/Q _6455_/B _6482_/A _8727_/Q vssd1 vssd1 vccd1 vccd1 _6457_/B sky130_fd_sc_hd__or4bb_1
X_6386_ _5491_/X _6380_/X _6383_/X _6385_/Y vssd1 vssd1 vccd1 vccd1 _8714_/D sky130_fd_sc_hd__a31oi_1
X_5406_ _5408_/B _5406_/B vssd1 vssd1 vccd1 vccd1 _8701_/D sky130_fd_sc_hd__nor2_1
X_8125_ _8124_/A _8124_/B _8124_/C vssd1 vssd1 vccd1 vccd1 _8126_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5337_ _8685_/Q _8684_/Q vssd1 vssd1 vccd1 vccd1 _6535_/A sky130_fd_sc_hd__or2_1
XFILLER_87_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8056_ _8056_/A _8056_/B vssd1 vssd1 vccd1 vccd1 _8135_/A sky130_fd_sc_hd__and2_1
X_5268_ _4950_/X _5164_/X _5261_/X _5265_/X _5267_/X vssd1 vssd1 vccd1 vccd1 _5268_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_102_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7007_ _7118_/B _7006_/X _6854_/A _7282_/A vssd1 vssd1 vccd1 vccd1 _7412_/A sky130_fd_sc_hd__o31ai_4
XFILLER_68_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5199_ _5199_/A _5199_/B vssd1 vssd1 vccd1 vccd1 _5199_/Y sky130_fd_sc_hd__nand2_1
XFILLER_71_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8958_ _8958_/A _4443_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[7] sky130_fd_sc_hd__ebufn_8
X_7909_ _7908_/B _7908_/C _7903_/A vssd1 vssd1 vccd1 vccd1 _7910_/C sky130_fd_sc_hd__a21o_1
XFILLER_70_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8889_ _8889_/A _4367_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[8] sky130_fd_sc_hd__ebufn_8
XFILLER_24_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4570_ _7700_/A _5298_/A _4870_/A _4823_/A vssd1 vssd1 vccd1 vccd1 _4692_/C sky130_fd_sc_hd__or4_1
X_6240_ _6158_/A _6158_/B _6159_/A vssd1 vssd1 vccd1 vccd1 _6240_/Y sky130_fd_sc_hd__a21oi_1
X_6171_ _6171_/A _6171_/B vssd1 vssd1 vccd1 vccd1 _6252_/B sky130_fd_sc_hd__nand2_1
X_5122_ _5250_/B _5112_/X _5121_/X vssd1 vssd1 vccd1 vccd1 _5122_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_69_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5053_ _5172_/A _5053_/B vssd1 vssd1 vccd1 vccd1 _5124_/D sky130_fd_sc_hd__nand2_1
XFILLER_84_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5955_ _5955_/A _5955_/B vssd1 vssd1 vccd1 vccd1 _5956_/B sky130_fd_sc_hd__xnor2_1
X_8743_ _8753_/CLK _8743_/D vssd1 vssd1 vccd1 vccd1 _8743_/Q sky130_fd_sc_hd__dfxtp_1
X_5886_ _5886_/A _5867_/X vssd1 vssd1 vccd1 vccd1 _5969_/B sky130_fd_sc_hd__or2b_1
X_8674_ _8785_/CLK _8674_/D vssd1 vssd1 vccd1 vccd1 _8674_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4906_ _5085_/A _5288_/B _5141_/C vssd1 vssd1 vccd1 vccd1 _5179_/B sky130_fd_sc_hd__or3b_4
XFILLER_33_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7625_ _8768_/Q _7649_/B _7624_/X vssd1 vssd1 vccd1 vccd1 _7625_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_21_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4837_ _4883_/B _4925_/B vssd1 vssd1 vccd1 vccd1 _5155_/C sky130_fd_sc_hd__nor2_2
X_7556_ _7556_/A _8746_/Q vssd1 vssd1 vccd1 vccd1 _7558_/B sky130_fd_sc_hd__xor2_1
X_4768_ _4765_/X _7576_/B _4768_/C vssd1 vssd1 vccd1 vccd1 _4769_/A sky130_fd_sc_hd__and3b_1
XFILLER_4_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7487_ _7487_/A _7487_/B vssd1 vssd1 vccd1 vccd1 _7487_/Y sky130_fd_sc_hd__nor2_1
X_6507_ _6506_/B _8737_/Q _6501_/B _8739_/Q vssd1 vssd1 vccd1 vccd1 _6508_/C sky130_fd_sc_hd__a31o_1
X_4699_ _5275_/A vssd1 vssd1 vccd1 vccd1 _5047_/A sky130_fd_sc_hd__clkbuf_2
X_6438_ _8741_/Q vssd1 vssd1 vccd1 vccd1 _6515_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_8874__91 vssd1 vssd1 vccd1 vccd1 _8874__91/HI _8983_/A sky130_fd_sc_hd__conb_1
X_6369_ _6369_/A _6369_/B _6369_/C vssd1 vssd1 vccd1 vccd1 _6369_/X sky130_fd_sc_hd__and3_1
X_8108_ _8420_/A vssd1 vssd1 vccd1 vccd1 _8236_/C sky130_fd_sc_hd__inv_2
XFILLER_88_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8039_ _8058_/A _8039_/B _8039_/C vssd1 vssd1 vccd1 vccd1 _8039_/X sky130_fd_sc_hd__or3_1
XFILLER_29_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5740_ _5620_/A _5619_/B _5620_/B _5739_/Y _5687_/A vssd1 vssd1 vccd1 vccd1 _5751_/A
+ sky130_fd_sc_hd__o311a_2
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5671_ _5799_/A _5671_/B vssd1 vssd1 vccd1 vccd1 _5673_/B sky130_fd_sc_hd__nand2_1
X_7410_ _7410_/A _7410_/B vssd1 vssd1 vccd1 vccd1 _7423_/A sky130_fd_sc_hd__xor2_1
X_8390_ _8461_/S _8390_/B vssd1 vssd1 vccd1 vccd1 _8463_/C sky130_fd_sc_hd__xnor2_2
X_4622_ _8632_/Q _8631_/Q _8633_/Q vssd1 vssd1 vccd1 vccd1 _4631_/C sky130_fd_sc_hd__and3_1
X_4553_ _7739_/B vssd1 vssd1 vccd1 vccd1 _4733_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_7341_ _7341_/A _7352_/A vssd1 vssd1 vccd1 vccd1 _7342_/B sky130_fd_sc_hd__xnor2_4
X_4484_ _4486_/A vssd1 vssd1 vccd1 vccd1 _4484_/Y sky130_fd_sc_hd__inv_2
X_7272_ _7272_/A _7409_/B _7272_/C vssd1 vssd1 vccd1 vccd1 _7276_/A sky130_fd_sc_hd__nand3_1
XFILLER_89_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6223_ _6177_/A _6177_/B _6178_/B _6178_/A vssd1 vssd1 vccd1 vccd1 _6343_/B sky130_fd_sc_hd__a2bb2o_1
X_6154_ _6154_/A _6154_/B vssd1 vssd1 vccd1 vccd1 _6235_/A sky130_fd_sc_hd__xnor2_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6085_ _6085_/A _6085_/B vssd1 vssd1 vccd1 vccd1 _6181_/B sky130_fd_sc_hd__xnor2_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5105_ _5176_/A vssd1 vssd1 vccd1 vccd1 _5150_/A sky130_fd_sc_hd__clkbuf_2
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5036_ _5036_/A _5036_/B _5238_/C vssd1 vssd1 vccd1 vccd1 _5038_/A sky130_fd_sc_hd__or3_2
XFILLER_72_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6987_ _7228_/A _6834_/B _6814_/B _6814_/A vssd1 vssd1 vccd1 vccd1 _7069_/A sky130_fd_sc_hd__a22o_1
XFILLER_41_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5938_ _5938_/A _5938_/B vssd1 vssd1 vccd1 vccd1 _5939_/B sky130_fd_sc_hd__nand2_1
XFILLER_13_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8726_ _8742_/CLK _8726_/D vssd1 vssd1 vccd1 vccd1 _8726_/Q sky130_fd_sc_hd__dfxtp_1
X_5869_ _5810_/X _5792_/X _5867_/X _5868_/Y vssd1 vssd1 vccd1 vccd1 _5885_/A sky130_fd_sc_hd__o211ai_2
X_8657_ _8778_/CLK _8657_/D vssd1 vssd1 vccd1 vccd1 _8657_/Q sky130_fd_sc_hd__dfxtp_2
X_7608_ _8769_/Q vssd1 vssd1 vccd1 vccd1 _7630_/A sky130_fd_sc_hd__clkbuf_2
X_8588_ _8588_/A _8778_/Q vssd1 vssd1 vccd1 vccd1 _8588_/Y sky130_fd_sc_hd__nor2_1
XFILLER_5_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7539_ _7539_/A _7551_/A _7539_/C vssd1 vssd1 vccd1 vccd1 _7539_/X sky130_fd_sc_hd__and3_1
XFILLER_0_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_9_0_wb_clk_i clkbuf_4_9_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _8784_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_79_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7890_ _7890_/A vssd1 vssd1 vccd1 vccd1 _8582_/A sky130_fd_sc_hd__inv_2
XFILLER_54_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6910_ _6910_/A _6910_/B _6910_/C vssd1 vssd1 vccd1 vccd1 _6910_/X sky130_fd_sc_hd__and3_1
XFILLER_47_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6841_ _6839_/X _6788_/B _6840_/X vssd1 vssd1 vccd1 vccd1 _6881_/B sky130_fd_sc_hd__a21o_1
X_8511_ _8279_/A _8393_/A _8465_/A vssd1 vssd1 vccd1 vccd1 _8512_/B sky130_fd_sc_hd__o21ba_1
X_6772_ _7123_/A _7020_/A vssd1 vssd1 vccd1 vccd1 _6965_/A sky130_fd_sc_hd__nand2_2
X_5723_ _6004_/A _5824_/B _5611_/B _5722_/Y vssd1 vssd1 vccd1 vccd1 _5730_/A sky130_fd_sc_hd__a31o_1
X_8442_ _8443_/A _8443_/B _8441_/Y vssd1 vssd1 vccd1 vccd1 _8442_/X sky130_fd_sc_hd__o21ba_1
X_5654_ _5700_/A _5916_/B vssd1 vssd1 vccd1 vccd1 _5666_/A sky130_fd_sc_hd__nand2_1
X_8373_ _8373_/A _8439_/C vssd1 vssd1 vccd1 vccd1 _8399_/A sky130_fd_sc_hd__xnor2_2
X_4605_ _8642_/Q _8641_/Q _8644_/Q _8643_/Q vssd1 vssd1 vccd1 vccd1 _4606_/D sky130_fd_sc_hd__or4_1
XFILLER_30_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5585_ _5585_/A _5585_/B vssd1 vssd1 vccd1 vccd1 _5688_/A sky130_fd_sc_hd__xnor2_4
X_7324_ _7484_/S _7237_/B _7323_/X vssd1 vssd1 vccd1 vccd1 _7341_/A sky130_fd_sc_hd__a21bo_2
X_4536_ _8665_/Q vssd1 vssd1 vccd1 vccd1 _6621_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_104_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4467_ _4468_/A vssd1 vssd1 vccd1 vccd1 _4467_/Y sky130_fd_sc_hd__inv_2
X_7255_ _7255_/A _7238_/A vssd1 vssd1 vccd1 vccd1 _7257_/A sky130_fd_sc_hd__or2b_1
XFILLER_104_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4398_ _4400_/A vssd1 vssd1 vccd1 vccd1 _4398_/Y sky130_fd_sc_hd__inv_2
X_6206_ _6207_/A _6207_/B _6207_/C vssd1 vssd1 vccd1 vccd1 _6208_/A sky130_fd_sc_hd__a21oi_1
X_8844__61 vssd1 vssd1 vccd1 vccd1 _8844__61/HI _8953_/A sky130_fd_sc_hd__conb_1
X_7186_ _7009_/S _7186_/B _7198_/A vssd1 vssd1 vccd1 vccd1 _7186_/X sky130_fd_sc_hd__and3b_1
X_6137_ _6137_/A _6137_/B vssd1 vssd1 vccd1 vccd1 _6137_/Y sky130_fd_sc_hd__nor2_1
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6068_ _6068_/A _6068_/B _6068_/C vssd1 vssd1 vccd1 vccd1 _6075_/A sky130_fd_sc_hd__and3_1
X_5019_ _5182_/A vssd1 vssd1 vccd1 vccd1 _5192_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_41_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8709_ _8783_/CLK _8709_/D vssd1 vssd1 vccd1 vccd1 _8709_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5370_ _8690_/Q _5372_/C _5360_/X vssd1 vssd1 vccd1 vccd1 _5371_/B sky130_fd_sc_hd__o21ai_1
XFILLER_99_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7040_ _7212_/A _7040_/B vssd1 vssd1 vccd1 vccd1 _7041_/B sky130_fd_sc_hd__xnor2_1
XFILLER_101_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7942_ _8325_/A _8348_/A vssd1 vssd1 vccd1 vccd1 _7955_/A sky130_fd_sc_hd__or2_1
XFILLER_70_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7873_ _8138_/A _7873_/B vssd1 vssd1 vccd1 vccd1 _8586_/A sky130_fd_sc_hd__nand2_1
X_6824_ _6891_/A _6891_/B _6823_/Y vssd1 vssd1 vccd1 vccd1 _6956_/A sky130_fd_sc_hd__o21ai_1
XFILLER_23_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6755_ _6755_/A _6755_/B vssd1 vssd1 vccd1 vccd1 _6755_/X sky130_fd_sc_hd__or2_1
X_5706_ _5710_/A _5710_/B vssd1 vssd1 vccd1 vccd1 _5711_/A sky130_fd_sc_hd__nand2_1
X_8425_ _8338_/B _8425_/B vssd1 vssd1 vccd1 vccd1 _8425_/X sky130_fd_sc_hd__and2b_1
X_6686_ _6858_/B vssd1 vssd1 vccd1 vccd1 _6834_/B sky130_fd_sc_hd__clkbuf_2
X_5637_ _5637_/A vssd1 vssd1 vccd1 vccd1 _6193_/A sky130_fd_sc_hd__clkbuf_2
X_8356_ _8358_/B _8356_/B vssd1 vssd1 vccd1 vccd1 _8420_/B sky130_fd_sc_hd__and2_1
X_5568_ _8719_/Q _7729_/B vssd1 vssd1 vccd1 vccd1 _5568_/X sky130_fd_sc_hd__and2b_1
X_8287_ _8320_/A _8320_/B vssd1 vssd1 vccd1 vccd1 _8306_/A sky130_fd_sc_hd__xor2_2
X_7307_ _7208_/A _7208_/B _7306_/X vssd1 vssd1 vccd1 vccd1 _7397_/B sky130_fd_sc_hd__o21bai_1
X_4519_ _5298_/A vssd1 vssd1 vccd1 vccd1 _4804_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5499_ _5552_/A _5526_/B _5498_/X vssd1 vssd1 vccd1 vccd1 _5547_/A sky130_fd_sc_hd__a21o_1
X_7238_ _7238_/A _7255_/A vssd1 vssd1 vccd1 vccd1 _7239_/B sky130_fd_sc_hd__xnor2_1
X_7169_ _7169_/A _7016_/B vssd1 vssd1 vccd1 vccd1 _7169_/X sky130_fd_sc_hd__or2b_1
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4870_ _4870_/A _4874_/A _4874_/B _4902_/C vssd1 vssd1 vccd1 vccd1 _4892_/A sky130_fd_sc_hd__or4b_1
XFILLER_20_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6540_ _8746_/Q vssd1 vssd1 vccd1 vccd1 _7578_/B sky130_fd_sc_hd__inv_2
X_6471_ _6471_/A vssd1 vssd1 vccd1 vccd1 _8727_/D sky130_fd_sc_hd__clkbuf_1
X_8210_ _8028_/A _8336_/A _8096_/B _8236_/A vssd1 vssd1 vccd1 vccd1 _8288_/B sky130_fd_sc_hd__a2bb2o_1
X_5422_ _6409_/A _6405_/A _8718_/Q _5421_/Y vssd1 vssd1 vccd1 vccd1 _5422_/X sky130_fd_sc_hd__a31o_1
X_8141_ _8054_/Y _8556_/B _8559_/B _8559_/A _8559_/C vssd1 vssd1 vccd1 vccd1 _8562_/B
+ sky130_fd_sc_hd__o2111ai_2
X_5353_ _5353_/A vssd1 vssd1 vccd1 vccd1 _8685_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8072_ _8008_/A _8258_/A _8011_/B _8157_/A vssd1 vssd1 vccd1 vccd1 _8078_/A sky130_fd_sc_hd__a22o_1
XFILLER_59_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5284_ _5077_/B _5077_/C _5283_/X _5087_/B _5215_/A vssd1 vssd1 vccd1 vccd1 _5285_/D
+ sky130_fd_sc_hd__o32a_1
X_8814__31 vssd1 vssd1 vccd1 vccd1 _8814__31/HI _8909_/A sky130_fd_sc_hd__conb_1
XFILLER_87_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_8 _5252_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7023_ _7023_/A _7023_/B vssd1 vssd1 vccd1 vccd1 _7024_/B sky130_fd_sc_hd__xnor2_2
XFILLER_67_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8974_ _8974_/A _4468_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[23] sky130_fd_sc_hd__ebufn_8
XFILLER_43_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7925_ _7925_/A vssd1 vssd1 vccd1 vccd1 _8376_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_82_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7856_ _7938_/A _7856_/B vssd1 vssd1 vccd1 vccd1 _7858_/A sky130_fd_sc_hd__and2b_1
XFILLER_51_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6807_ _6807_/A _6807_/B vssd1 vssd1 vccd1 vccd1 _6807_/X sky130_fd_sc_hd__and2_1
X_7787_ _8450_/A _7924_/A vssd1 vssd1 vccd1 vccd1 _7820_/A sky130_fd_sc_hd__nand2_1
X_4999_ _5136_/C vssd1 vssd1 vccd1 vccd1 _5224_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6738_ _6632_/A _6632_/B _6764_/B _6737_/X vssd1 vssd1 vccd1 vccd1 _6775_/B sky130_fd_sc_hd__a31o_4
X_6669_ _6886_/A vssd1 vssd1 vccd1 vccd1 _6814_/A sky130_fd_sc_hd__clkbuf_2
X_8408_ _8405_/A _8408_/B vssd1 vssd1 vccd1 vccd1 _8477_/B sky130_fd_sc_hd__and2b_1
X_8339_ _8339_/A _8339_/B vssd1 vssd1 vccd1 vccd1 _8341_/A sky130_fd_sc_hd__nand2_1
XFILLER_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5971_ _5971_/A _5971_/B vssd1 vssd1 vccd1 vccd1 _5971_/Y sky130_fd_sc_hd__nand2_1
XFILLER_92_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7710_ _7946_/A _8325_/B _8354_/A _7854_/A vssd1 vssd1 vccd1 vccd1 _7710_/X sky130_fd_sc_hd__or4b_2
XFILLER_52_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8690_ _8704_/CLK _8690_/D vssd1 vssd1 vccd1 vccd1 _8690_/Q sky130_fd_sc_hd__dfxtp_1
X_4922_ _4922_/A _4935_/B vssd1 vssd1 vccd1 vccd1 _5077_/C sky130_fd_sc_hd__nor2_2
X_7641_ _8603_/A _7641_/B vssd1 vssd1 vccd1 vccd1 _7641_/X sky130_fd_sc_hd__or2_1
XFILLER_100_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4853_ _4937_/B vssd1 vssd1 vccd1 vccd1 _5050_/D sky130_fd_sc_hd__clkbuf_2
X_4784_ _4784_/A vssd1 vssd1 vccd1 vccd1 _5040_/A sky130_fd_sc_hd__buf_2
X_7572_ _6660_/A _8746_/Q _7569_/B vssd1 vssd1 vccd1 vccd1 _7572_/X sky130_fd_sc_hd__o21a_1
X_6523_ _8744_/Q _6521_/A _6522_/Y _5335_/X vssd1 vssd1 vccd1 vccd1 _8744_/D sky130_fd_sc_hd__o211a_1
X_6454_ _8730_/Q _8736_/Q _6454_/C _6454_/D vssd1 vssd1 vccd1 vccd1 _7619_/B sky130_fd_sc_hd__or4_4
X_5405_ _8701_/Q _5404_/B _5392_/X vssd1 vssd1 vccd1 vccd1 _5406_/B sky130_fd_sc_hd__o21ai_1
X_6385_ _8574_/A _8714_/Q vssd1 vssd1 vccd1 vccd1 _6385_/Y sky130_fd_sc_hd__nor2_1
X_8124_ _8124_/A _8124_/B _8124_/C vssd1 vssd1 vccd1 vccd1 _8304_/A sky130_fd_sc_hd__and3_1
X_5336_ _8758_/Q _5320_/A _5334_/X _5335_/X vssd1 vssd1 vccd1 vccd1 _8683_/D sky130_fd_sc_hd__o211a_1
X_8055_ _8055_/A _8053_/B vssd1 vssd1 vccd1 vccd1 _8311_/A sky130_fd_sc_hd__or2b_1
X_5267_ _5266_/A _5261_/B _5171_/B _5266_/Y vssd1 vssd1 vccd1 vccd1 _5267_/X sky130_fd_sc_hd__o31a_1
X_7006_ _7279_/A vssd1 vssd1 vccd1 vccd1 _7006_/X sky130_fd_sc_hd__clkbuf_2
X_5198_ _5280_/A _5288_/C vssd1 vssd1 vccd1 vccd1 _5199_/B sky130_fd_sc_hd__nor2_1
XFILLER_83_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8957_ _8957_/A _4441_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[6] sky130_fd_sc_hd__ebufn_8
XFILLER_83_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7908_ _8008_/A _7908_/B _7908_/C vssd1 vssd1 vccd1 vccd1 _7910_/B sky130_fd_sc_hd__nand3_1
XFILLER_55_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8888_ _8888_/A _4366_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[7] sky130_fd_sc_hd__ebufn_8
XFILLER_24_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7839_ _7854_/A _7839_/B _7854_/B vssd1 vssd1 vccd1 vccd1 _7839_/X sky130_fd_sc_hd__and3_1
XFILLER_34_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_4_11_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8771_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6170_ _6172_/A vssd1 vssd1 vccd1 vccd1 _6251_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_69_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5121_ _5116_/X _5120_/X _4733_/C _5135_/A _5059_/B vssd1 vssd1 vccd1 vccd1 _5121_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_97_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5052_ _5088_/B _5066_/B vssd1 vssd1 vccd1 vccd1 _5277_/B sky130_fd_sc_hd__nand2_1
XFILLER_92_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8742_ _8742_/CLK _8742_/D vssd1 vssd1 vccd1 vccd1 _8742_/Q sky130_fd_sc_hd__dfxtp_1
X_5954_ _6047_/A _5954_/B vssd1 vssd1 vccd1 vccd1 _5955_/B sky130_fd_sc_hd__nor2_1
XFILLER_52_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5885_ _5885_/A _5885_/B vssd1 vssd1 vccd1 vccd1 _5967_/B sky130_fd_sc_hd__nand2_1
XFILLER_80_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8673_ _8785_/CLK _8673_/D vssd1 vssd1 vccd1 vccd1 _8673_/Q sky130_fd_sc_hd__dfxtp_1
X_4905_ _5288_/C _5088_/A vssd1 vssd1 vccd1 vccd1 _5141_/C sky130_fd_sc_hd__and2b_1
XFILLER_21_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7624_ _7656_/B vssd1 vssd1 vccd1 vccd1 _7624_/X sky130_fd_sc_hd__clkbuf_2
X_4836_ _4836_/A vssd1 vssd1 vccd1 vccd1 _4883_/B sky130_fd_sc_hd__buf_2
X_7555_ _7555_/A vssd1 vssd1 vccd1 vccd1 _8759_/D sky130_fd_sc_hd__clkbuf_1
X_6506_ _8739_/Q _6506_/B _6506_/C vssd1 vssd1 vccd1 vccd1 _6510_/B sky130_fd_sc_hd__and3_1
X_4767_ _5100_/A _4767_/B vssd1 vssd1 vccd1 vccd1 _4768_/C sky130_fd_sc_hd__or2_1
X_7486_ _7486_/A _7486_/B vssd1 vssd1 vccd1 vccd1 _7502_/A sky130_fd_sc_hd__xnor2_1
X_4698_ _8653_/Q vssd1 vssd1 vccd1 vccd1 _5210_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6437_ _8725_/Q vssd1 vssd1 vccd1 vccd1 _6455_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6368_ _6369_/B _6369_/C _6369_/A vssd1 vssd1 vccd1 vccd1 _6368_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_88_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8107_ _8121_/B _8124_/B vssd1 vssd1 vccd1 vccd1 _8110_/A sky130_fd_sc_hd__or2b_1
X_5319_ _8775_/Q _5307_/X _5318_/X _5311_/X vssd1 vssd1 vccd1 vccd1 _8676_/D sky130_fd_sc_hd__o211a_1
X_6299_ _6292_/A _6297_/A _6292_/B vssd1 vssd1 vccd1 vccd1 _6358_/B sky130_fd_sc_hd__a21bo_1
XFILLER_29_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8038_ _8119_/A _8038_/B vssd1 vssd1 vccd1 vccd1 _8039_/C sky130_fd_sc_hd__xor2_1
XFILLER_29_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5670_ _5670_/A _5670_/B vssd1 vssd1 vccd1 vccd1 _5671_/B sky130_fd_sc_hd__nand2_1
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4621_ _4621_/A vssd1 vssd1 vccd1 vccd1 _8632_/D sky130_fd_sc_hd__clkbuf_1
X_4552_ _8655_/Q vssd1 vssd1 vccd1 vccd1 _7739_/B sky130_fd_sc_hd__buf_4
X_7340_ _7340_/A _7340_/B vssd1 vssd1 vccd1 vccd1 _7352_/A sky130_fd_sc_hd__xnor2_2
X_4483_ _4486_/A vssd1 vssd1 vccd1 vccd1 _4483_/Y sky130_fd_sc_hd__inv_2
X_7271_ _7409_/A _7270_/C _7261_/A vssd1 vssd1 vccd1 vccd1 _7272_/C sky130_fd_sc_hd__a21o_1
X_6222_ _6213_/A _6213_/B _6221_/X vssd1 vssd1 vccd1 vccd1 _6351_/A sky130_fd_sc_hd__a21o_1
XFILLER_97_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6153_ _6171_/A _6153_/B vssd1 vssd1 vccd1 vccd1 _6154_/B sky130_fd_sc_hd__xnor2_1
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6084_ _6092_/A _6194_/A vssd1 vssd1 vccd1 vccd1 _6085_/B sky130_fd_sc_hd__xor2_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5104_ _5231_/A _5228_/B _5093_/X _5103_/X _4819_/A vssd1 vssd1 vccd1 vccd1 _5130_/C
+ sky130_fd_sc_hd__o311a_1
XFILLER_85_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5035_ _5206_/A _5211_/A vssd1 vssd1 vccd1 vccd1 _5238_/C sky130_fd_sc_hd__or2_1
XFILLER_38_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6986_ _6988_/B _6988_/A vssd1 vssd1 vccd1 vccd1 _7067_/B sky130_fd_sc_hd__or2b_1
XFILLER_25_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5937_ _5937_/A _5937_/B vssd1 vssd1 vccd1 vccd1 _5938_/B sky130_fd_sc_hd__or2_1
X_8725_ _8742_/CLK _8725_/D vssd1 vssd1 vccd1 vccd1 _8725_/Q sky130_fd_sc_hd__dfxtp_1
X_8656_ _8778_/CLK _8656_/D vssd1 vssd1 vccd1 vccd1 _8656_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_15_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5868_ _5886_/A _5867_/B _5867_/C vssd1 vssd1 vccd1 vccd1 _5868_/Y sky130_fd_sc_hd__o21ai_1
X_7607_ _8773_/Q vssd1 vssd1 vccd1 vccd1 _7775_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5799_ _5799_/A _5799_/B vssd1 vssd1 vccd1 vccd1 _5800_/B sky130_fd_sc_hd__nand2_1
X_8587_ _7887_/Y _8586_/B _8586_/Y _8578_/A _8578_/B vssd1 vssd1 vccd1 vccd1 _8587_/X
+ sky130_fd_sc_hd__a2111o_1
X_4819_ _4819_/A vssd1 vssd1 vccd1 vccd1 _4819_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_5_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7538_ _7538_/A _7544_/B vssd1 vssd1 vccd1 vccd1 _7539_/C sky130_fd_sc_hd__nand2_1
X_7469_ _7469_/A _7469_/B vssd1 vssd1 vccd1 vccd1 _7470_/B sky130_fd_sc_hd__xnor2_1
XFILLER_88_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6840_ _6840_/A _6840_/B vssd1 vssd1 vccd1 vccd1 _6840_/X sky130_fd_sc_hd__and2_1
XFILLER_35_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6771_ _6866_/C vssd1 vssd1 vccd1 vccd1 _7020_/A sky130_fd_sc_hd__clkbuf_2
X_8510_ _8510_/A _8510_/B vssd1 vssd1 vccd1 vccd1 _8537_/A sky130_fd_sc_hd__xnor2_1
X_5722_ _6263_/A _5984_/C vssd1 vssd1 vccd1 vccd1 _5722_/Y sky130_fd_sc_hd__nor2_1
X_8441_ _8441_/A _8527_/B vssd1 vssd1 vccd1 vccd1 _8441_/Y sky130_fd_sc_hd__xnor2_1
X_5653_ _5925_/B vssd1 vssd1 vccd1 vccd1 _5916_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8372_ _8438_/B _8372_/B vssd1 vssd1 vccd1 vccd1 _8439_/C sky130_fd_sc_hd__xnor2_1
X_5584_ _5680_/A _5584_/B vssd1 vssd1 vccd1 vccd1 _6378_/C sky130_fd_sc_hd__and2_2
X_4604_ _8651_/Q vssd1 vssd1 vccd1 vccd1 _5462_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_7_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7323_ _7323_/A _7236_/A vssd1 vssd1 vccd1 vccd1 _7323_/X sky130_fd_sc_hd__or2b_1
X_4535_ _4872_/B _4762_/A vssd1 vssd1 vccd1 vccd1 _4850_/A sky130_fd_sc_hd__and2_1
X_4466_ _4468_/A vssd1 vssd1 vccd1 vccd1 _4466_/Y sky130_fd_sc_hd__inv_2
X_7254_ _7242_/A _7242_/B _7253_/X vssd1 vssd1 vccd1 vccd1 _7345_/A sky130_fd_sc_hd__a21boi_1
X_4397_ _4400_/A vssd1 vssd1 vccd1 vccd1 _4397_/Y sky130_fd_sc_hd__inv_2
X_6205_ _6205_/A _6205_/B vssd1 vssd1 vccd1 vccd1 _6207_/C sky130_fd_sc_hd__xnor2_1
X_7185_ _7185_/A _7274_/A vssd1 vssd1 vccd1 vccd1 _7190_/A sky130_fd_sc_hd__xor2_1
X_6136_ _6120_/B _6122_/B _6120_/A vssd1 vssd1 vccd1 vccd1 _6215_/A sky130_fd_sc_hd__o21ba_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6067_ _6009_/A _6009_/B _6066_/X vssd1 vssd1 vccd1 vccd1 _6103_/A sky130_fd_sc_hd__a21oi_2
XFILLER_58_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5018_ _5163_/B _5014_/X _5017_/X _4967_/X vssd1 vssd1 vccd1 vccd1 _5018_/X sky130_fd_sc_hd__o22a_1
XFILLER_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6969_ _6967_/A _6967_/B _6975_/A vssd1 vssd1 vccd1 vccd1 _6971_/A sky130_fd_sc_hd__a21bo_1
XFILLER_41_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8708_ _8783_/CLK _8708_/D vssd1 vssd1 vccd1 vccd1 _8708_/Q sky130_fd_sc_hd__dfxtp_2
X_8639_ _8730_/CLK _8639_/D vssd1 vssd1 vccd1 vccd1 _8639_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7941_ _7854_/B _7850_/B _7940_/X vssd1 vssd1 vccd1 vccd1 _7951_/A sky130_fd_sc_hd__a21oi_1
XFILLER_82_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7872_ _7872_/A _7872_/B _7875_/A vssd1 vssd1 vccd1 vccd1 _7873_/B sky130_fd_sc_hd__or3_1
XFILLER_23_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6823_ _6823_/A _6823_/B vssd1 vssd1 vccd1 vccd1 _6823_/Y sky130_fd_sc_hd__nand2_1
XFILLER_50_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6754_ _6755_/B _6732_/X vssd1 vssd1 vccd1 vccd1 _6775_/A sky130_fd_sc_hd__nor2b_4
X_5705_ _6377_/A _6377_/B _6381_/B vssd1 vssd1 vccd1 vccd1 _5710_/B sky130_fd_sc_hd__and3_1
XFILLER_50_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6685_ _6707_/A _7416_/A vssd1 vssd1 vccd1 vccd1 _6858_/B sky130_fd_sc_hd__nor2_1
X_8424_ _8424_/A _8424_/B vssd1 vssd1 vccd1 vccd1 _8427_/A sky130_fd_sc_hd__xnor2_1
X_5636_ _5819_/C _5819_/D vssd1 vssd1 vccd1 vccd1 _5637_/A sky130_fd_sc_hd__nor2_1
XFILLER_12_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8355_ _8355_/A _8355_/B vssd1 vssd1 vccd1 vccd1 _8356_/B sky130_fd_sc_hd__nand2_1
X_5567_ _8719_/Q _7729_/B vssd1 vssd1 vccd1 vccd1 _5680_/B sky130_fd_sc_hd__xnor2_4
X_8286_ _8286_/A _8286_/B vssd1 vssd1 vccd1 vccd1 _8320_/B sky130_fd_sc_hd__xnor2_2
X_5498_ _8708_/Q _6630_/B vssd1 vssd1 vccd1 vccd1 _5498_/X sky130_fd_sc_hd__and2b_1
XFILLER_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7306_ _7382_/A _7306_/B vssd1 vssd1 vccd1 vccd1 _7306_/X sky130_fd_sc_hd__and2_1
X_4518_ _4902_/C vssd1 vssd1 vccd1 vccd1 _5298_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4449_ _4450_/A vssd1 vssd1 vccd1 vccd1 _4449_/Y sky130_fd_sc_hd__inv_2
X_7237_ _7484_/S _7237_/B vssd1 vssd1 vccd1 vccd1 _7255_/A sky130_fd_sc_hd__xnor2_1
X_7168_ _7168_/A _7168_/B vssd1 vssd1 vccd1 vccd1 _7219_/B sky130_fd_sc_hd__nand2_1
X_6119_ _6119_/A _6119_/B _6119_/C vssd1 vssd1 vccd1 vccd1 _6120_/B sky130_fd_sc_hd__nor3_1
XFILLER_85_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7099_ _7099_/A _7099_/B vssd1 vssd1 vccd1 vccd1 _7100_/B sky130_fd_sc_hd__and2_1
XFILLER_85_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6470_ _6473_/B _6470_/B _6508_/B vssd1 vssd1 vccd1 vccd1 _6471_/A sky130_fd_sc_hd__and3b_1
X_5421_ _6423_/A vssd1 vssd1 vccd1 vccd1 _5421_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8140_ _8138_/A _8139_/B _8556_/A _8137_/X vssd1 vssd1 vccd1 vccd1 _8559_/C sky130_fd_sc_hd__a2bb2o_1
X_5352_ _6535_/A _5409_/A _5352_/C vssd1 vssd1 vccd1 vccd1 _5353_/A sky130_fd_sc_hd__and3_1
X_8071_ _8151_/A _8151_/B vssd1 vssd1 vccd1 vccd1 _8080_/A sky130_fd_sc_hd__xnor2_1
XFILLER_101_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7022_ _7022_/A _7198_/C vssd1 vssd1 vccd1 vccd1 _7023_/B sky130_fd_sc_hd__xnor2_1
X_5283_ _5283_/A _5283_/B _5283_/C vssd1 vssd1 vccd1 vccd1 _5283_/X sky130_fd_sc_hd__or3_1
XFILLER_99_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_9 _6621_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8973_ _8973_/A _4467_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[22] sky130_fd_sc_hd__ebufn_8
XFILLER_55_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7924_ _7924_/A _8158_/A _7924_/C vssd1 vssd1 vccd1 vccd1 _7928_/B sky130_fd_sc_hd__and3_1
XFILLER_55_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7855_ _7940_/C _7855_/B vssd1 vssd1 vccd1 vccd1 _7856_/B sky130_fd_sc_hd__xor2_1
XFILLER_70_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6806_ _6807_/A _6807_/B vssd1 vssd1 vccd1 vccd1 _6845_/B sky130_fd_sc_hd__xor2_2
X_7786_ _8155_/A vssd1 vssd1 vccd1 vccd1 _8450_/A sky130_fd_sc_hd__clkbuf_2
X_4998_ _5272_/C vssd1 vssd1 vccd1 vccd1 _5136_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_23_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6737_ _6577_/A _7679_/A _6736_/X _6735_/B vssd1 vssd1 vccd1 vccd1 _6737_/X sky130_fd_sc_hd__a31o_1
X_6668_ _6799_/A vssd1 vssd1 vccd1 vccd1 _6886_/A sky130_fd_sc_hd__clkbuf_2
X_8407_ _8404_/B _8407_/B vssd1 vssd1 vccd1 vccd1 _8477_/A sky130_fd_sc_hd__and2b_1
X_5619_ _5619_/A _5619_/B vssd1 vssd1 vccd1 vccd1 _5634_/B sky130_fd_sc_hd__nor2_1
X_6599_ _6599_/A _6598_/X vssd1 vssd1 vccd1 vccd1 _6599_/X sky130_fd_sc_hd__or2b_1
X_8338_ _8425_/B _8338_/B vssd1 vssd1 vccd1 vccd1 _8342_/A sky130_fd_sc_hd__xor2_1
X_8269_ _8268_/B _8268_/C _8268_/A vssd1 vssd1 vccd1 vccd1 _8280_/B sky130_fd_sc_hd__a21o_1
XFILLER_78_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5970_ _5955_/A _5955_/B _5969_/X vssd1 vssd1 vccd1 vccd1 _6050_/A sky130_fd_sc_hd__a21oi_1
XFILLER_64_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4921_ _4921_/A _4925_/B vssd1 vssd1 vccd1 vccd1 _5148_/B sky130_fd_sc_hd__nor2_2
X_7640_ _7652_/C _7640_/B vssd1 vssd1 vccd1 vccd1 _7641_/B sky130_fd_sc_hd__xnor2_1
X_4852_ _4910_/B _4925_/B vssd1 vssd1 vccd1 vccd1 _4937_/B sky130_fd_sc_hd__nor2_1
XFILLER_45_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4783_ _4877_/C _4812_/B vssd1 vssd1 vccd1 vccd1 _4784_/A sky130_fd_sc_hd__or2_2
X_7571_ _7585_/A _7579_/B vssd1 vssd1 vccd1 vccd1 _7575_/A sky130_fd_sc_hd__xnor2_1
X_6522_ _8744_/Q _6521_/A _8745_/Q vssd1 vssd1 vccd1 vccd1 _6522_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6453_ _8734_/Q _8738_/Q _8737_/Q _8733_/Q vssd1 vssd1 vccd1 vccd1 _6454_/D sky130_fd_sc_hd__or4bb_1
X_5404_ _8701_/Q _5404_/B vssd1 vssd1 vccd1 vccd1 _5408_/B sky130_fd_sc_hd__and2_1
X_8123_ _8099_/A _8034_/A _8122_/Y vssd1 vssd1 vccd1 vccd1 _8124_/C sky130_fd_sc_hd__o21a_1
X_6384_ _7656_/B vssd1 vssd1 vccd1 vccd1 _8574_/A sky130_fd_sc_hd__clkbuf_2
X_5335_ _5335_/A vssd1 vssd1 vccd1 vccd1 _5335_/X sky130_fd_sc_hd__buf_2
X_8054_ _8556_/A vssd1 vssd1 vccd1 vccd1 _8054_/Y sky130_fd_sc_hd__inv_2
X_5266_ _5266_/A _5266_/B vssd1 vssd1 vccd1 vccd1 _5266_/Y sky130_fd_sc_hd__nand2_1
XFILLER_75_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7005_ _7288_/A _7005_/B vssd1 vssd1 vccd1 vccd1 _7014_/A sky130_fd_sc_hd__nand2_1
XFILLER_68_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5197_ _5197_/A _5274_/B _5197_/C _5197_/D vssd1 vssd1 vccd1 vccd1 _5197_/X sky130_fd_sc_hd__or4_2
XFILLER_28_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8956_ _8956_/A _4438_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[5] sky130_fd_sc_hd__ebufn_8
XFILLER_43_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7907_ _8073_/A _7907_/B vssd1 vssd1 vccd1 vccd1 _7908_/C sky130_fd_sc_hd__nand2_1
XFILLER_70_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8887_ _8887_/A _4365_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[6] sky130_fd_sc_hd__ebufn_8
XFILLER_34_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7838_ _8330_/A _8354_/A vssd1 vssd1 vccd1 vccd1 _7854_/B sky130_fd_sc_hd__nor2_2
XFILLER_51_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7769_ _7934_/A _7880_/A _7836_/C _8165_/B vssd1 vssd1 vccd1 vccd1 _7882_/B sky130_fd_sc_hd__o211ai_2
XFILLER_7_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5120_ _5148_/B _5120_/B _5190_/C _5197_/C vssd1 vssd1 vccd1 vccd1 _5120_/X sky130_fd_sc_hd__or4_1
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5051_ _5159_/B _5174_/A _5126_/D _5051_/D vssd1 vssd1 vccd1 vccd1 _5051_/X sky130_fd_sc_hd__or4_1
XFILLER_65_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8741_ _8742_/CLK _8741_/D vssd1 vssd1 vccd1 vccd1 _8741_/Q sky130_fd_sc_hd__dfxtp_1
X_5953_ _5953_/A _5953_/B vssd1 vssd1 vccd1 vccd1 _5954_/B sky130_fd_sc_hd__and2_1
XFILLER_52_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5884_ _5884_/A _5884_/B vssd1 vssd1 vccd1 vccd1 _5957_/A sky130_fd_sc_hd__and2_1
X_8672_ _8776_/CLK _8672_/D vssd1 vssd1 vccd1 vccd1 _8672_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4904_ _5100_/B _5009_/C _5119_/A vssd1 vssd1 vccd1 vccd1 _5088_/A sky130_fd_sc_hd__a21oi_4
XFILLER_33_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7623_ _7649_/B vssd1 vssd1 vccd1 vccd1 _8609_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_21_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4835_ _7672_/B _8664_/Q _8663_/Q _8662_/Q vssd1 vssd1 vccd1 vccd1 _4836_/A sky130_fd_sc_hd__or4_1
XFILLER_21_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7554_ _6567_/A _6568_/A _7558_/A vssd1 vssd1 vccd1 vccd1 _7555_/A sky130_fd_sc_hd__mux2_1
X_4766_ _4807_/A vssd1 vssd1 vccd1 vccd1 _7576_/B sky130_fd_sc_hd__clkbuf_2
X_6505_ _6506_/B _6506_/C _6504_/Y vssd1 vssd1 vccd1 vccd1 _8738_/D sky130_fd_sc_hd__a21oi_1
X_7485_ _7485_/A _7485_/B vssd1 vssd1 vccd1 vccd1 _7486_/B sky130_fd_sc_hd__xnor2_1
XFILLER_20_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4697_ _5231_/A _4697_/B vssd1 vssd1 vccd1 vccd1 _4702_/C sky130_fd_sc_hd__nand2_1
X_6436_ _6436_/A vssd1 vssd1 vccd1 vccd1 _8724_/D sky130_fd_sc_hd__clkbuf_1
X_6367_ _6367_/A _6367_/B _6367_/C vssd1 vssd1 vccd1 vccd1 _6367_/X sky130_fd_sc_hd__and3_1
X_8106_ _8325_/B _8028_/A _8343_/A vssd1 vssd1 vccd1 vccd1 _8124_/B sky130_fd_sc_hd__a21o_1
X_5318_ _8676_/Q _5326_/B vssd1 vssd1 vccd1 vccd1 _5318_/X sky130_fd_sc_hd__or2_1
XFILLER_102_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6298_ _6360_/B _6360_/C _6361_/B _6360_/A vssd1 vssd1 vccd1 vccd1 _6358_/A sky130_fd_sc_hd__a211o_1
XFILLER_88_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8037_ _7958_/A _7958_/B _8036_/Y vssd1 vssd1 vccd1 vccd1 _8038_/B sky130_fd_sc_hd__o21ai_1
X_5249_ _5249_/A _5249_/B vssd1 vssd1 vccd1 vccd1 _5301_/C sky130_fd_sc_hd__nand2_1
XFILLER_102_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8939_ _8939_/A _4428_/Y vssd1 vssd1 vccd1 vccd1 io_out[26] sky130_fd_sc_hd__ebufn_8
XFILLER_45_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8865__82 vssd1 vssd1 vccd1 vccd1 _8865__82/HI _8974_/A sky130_fd_sc_hd__conb_1
XFILLER_79_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4620_ _4620_/A _4679_/A _4620_/C vssd1 vssd1 vccd1 vccd1 _4621_/A sky130_fd_sc_hd__and3_1
X_4551_ _5301_/A _4754_/A vssd1 vssd1 vccd1 vccd1 _4566_/A sky130_fd_sc_hd__or2_1
X_4482_ _4486_/A vssd1 vssd1 vccd1 vccd1 _4482_/Y sky130_fd_sc_hd__inv_2
X_7270_ _7405_/A _7409_/A _7270_/C vssd1 vssd1 vccd1 vccd1 _7409_/B sky130_fd_sc_hd__nand3_1
X_6221_ _6212_/A _6221_/B vssd1 vssd1 vccd1 vccd1 _6221_/X sky130_fd_sc_hd__and2b_1
X_6152_ _6152_/A _6152_/B vssd1 vssd1 vccd1 vccd1 _6154_/A sky130_fd_sc_hd__xor2_1
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5103_ _5095_/X _5102_/X _4720_/A vssd1 vssd1 vccd1 vccd1 _5103_/X sky130_fd_sc_hd__a21o_1
XFILLER_85_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6083_ _5625_/B _6274_/B _5981_/B _6068_/B vssd1 vssd1 vccd1 vccd1 _6181_/A sky130_fd_sc_hd__a22o_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5034_ _5179_/B _5228_/B vssd1 vssd1 vccd1 vccd1 _5036_/B sky130_fd_sc_hd__or2_1
XFILLER_25_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6985_ _7090_/A _7090_/B _6984_/X vssd1 vssd1 vccd1 vccd1 _6988_/A sky130_fd_sc_hd__a21bo_1
XFILLER_25_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5936_ _5936_/A _5936_/B vssd1 vssd1 vccd1 vccd1 _5938_/A sky130_fd_sc_hd__nand2_1
XFILLER_15_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8724_ _8730_/CLK _8724_/D vssd1 vssd1 vccd1 vccd1 _8724_/Q sky130_fd_sc_hd__dfxtp_1
X_8655_ _8778_/CLK _8655_/D vssd1 vssd1 vccd1 vccd1 _8655_/Q sky130_fd_sc_hd__dfxtp_2
X_5867_ _5886_/A _5867_/B _5867_/C vssd1 vssd1 vccd1 vccd1 _5867_/X sky130_fd_sc_hd__or3_1
X_7606_ _7606_/A _7606_/B _7606_/C vssd1 vssd1 vccd1 vccd1 _8766_/D sky130_fd_sc_hd__nand3_1
XFILLER_21_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5798_ _5799_/A _5799_/B vssd1 vssd1 vccd1 vccd1 _5879_/A sky130_fd_sc_hd__or2_1
X_8586_ _8586_/A _8586_/B vssd1 vssd1 vccd1 vccd1 _8586_/Y sky130_fd_sc_hd__nor2_1
X_4818_ _4818_/A _4818_/B vssd1 vssd1 vccd1 vccd1 _4819_/A sky130_fd_sc_hd__nor2_1
X_7537_ _7537_/A _7537_/B vssd1 vssd1 vccd1 vccd1 _7544_/B sky130_fd_sc_hd__nor2_1
X_4749_ _5249_/A vssd1 vssd1 vccd1 vccd1 _5300_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_7468_ _7309_/A _7388_/S _7389_/B _6813_/B vssd1 vssd1 vccd1 vccd1 _7469_/B sky130_fd_sc_hd__a22o_1
X_6419_ _8721_/Q _5462_/X _6418_/X _5335_/X vssd1 vssd1 vccd1 vccd1 _8721_/D sky130_fd_sc_hd__o211a_1
X_7399_ _7399_/A _7399_/B vssd1 vssd1 vccd1 vccd1 _7473_/A sky130_fd_sc_hd__xnor2_2
XFILLER_103_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6770_ _6770_/A _6770_/B vssd1 vssd1 vccd1 vccd1 _6866_/C sky130_fd_sc_hd__xnor2_2
X_5721_ _5627_/A _5627_/B _5720_/Y vssd1 vssd1 vccd1 vccd1 _5746_/A sky130_fd_sc_hd__a21bo_1
XFILLER_50_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8440_ _8496_/S _8356_/B _8358_/B vssd1 vssd1 vccd1 vccd1 _8527_/B sky130_fd_sc_hd__a21bo_1
X_5652_ _5769_/A _5652_/B vssd1 vssd1 vccd1 vccd1 _5925_/B sky130_fd_sc_hd__xnor2_1
X_8371_ _8371_/A _8371_/B vssd1 vssd1 vccd1 vccd1 _8372_/B sky130_fd_sc_hd__xnor2_1
X_5583_ _6004_/A vssd1 vssd1 vccd1 vccd1 _6378_/D sky130_fd_sc_hd__clkbuf_1
X_4603_ _4807_/A vssd1 vssd1 vccd1 vccd1 _4615_/A sky130_fd_sc_hd__buf_2
X_7322_ _7354_/B _7322_/B vssd1 vssd1 vccd1 vccd1 _7342_/A sky130_fd_sc_hd__xnor2_2
X_4534_ _4878_/C vssd1 vssd1 vccd1 vccd1 _4762_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_7_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4465_ _4468_/A vssd1 vssd1 vccd1 vccd1 _4465_/Y sky130_fd_sc_hd__inv_2
X_7253_ _7253_/A _7241_/A vssd1 vssd1 vccd1 vccd1 _7253_/X sky130_fd_sc_hd__or2b_1
X_4396_ _4400_/A vssd1 vssd1 vccd1 vccd1 _4396_/Y sky130_fd_sc_hd__inv_2
X_6204_ _6204_/A _6204_/B vssd1 vssd1 vccd1 vccd1 _6205_/B sky130_fd_sc_hd__nor2_1
X_7184_ _7288_/A _7288_/B vssd1 vssd1 vccd1 vccd1 _7192_/A sky130_fd_sc_hd__xor2_2
X_6135_ _6125_/A _6125_/B _6134_/Y vssd1 vssd1 vccd1 vccd1 _6294_/A sky130_fd_sc_hd__a21o_1
XFILLER_97_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6066_ _6001_/A _6066_/B vssd1 vssd1 vccd1 vccd1 _6066_/X sky130_fd_sc_hd__and2b_1
XFILLER_58_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5017_ _5047_/A _5157_/B _4987_/X _5174_/B vssd1 vssd1 vccd1 vccd1 _5017_/X sky130_fd_sc_hd__a211o_1
XFILLER_45_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8707_ _8720_/CLK _8707_/D vssd1 vssd1 vccd1 vccd1 _8707_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6968_ _7080_/D _6968_/B _6967_/X vssd1 vssd1 vccd1 vccd1 _6975_/A sky130_fd_sc_hd__or3b_1
X_5919_ _5856_/A _6171_/A _5918_/X vssd1 vssd1 vccd1 vccd1 _5920_/B sky130_fd_sc_hd__o21ba_1
X_6899_ _6757_/A _6757_/B _6757_/C _6851_/Y _6765_/A vssd1 vssd1 vccd1 vccd1 _6900_/A
+ sky130_fd_sc_hd__o311a_1
XFILLER_42_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8638_ _8730_/CLK _8638_/D vssd1 vssd1 vccd1 vccd1 _8638_/Q sky130_fd_sc_hd__dfxtp_1
X_8569_ _8571_/A _8567_/X _8568_/X vssd1 vssd1 vccd1 vccd1 _8576_/B sky130_fd_sc_hd__a21oi_1
X_8835__52 vssd1 vssd1 vccd1 vccd1 _8835__52/HI _8944_/A sky130_fd_sc_hd__conb_1
XFILLER_88_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7940_ _7940_/A _8098_/A _7940_/C vssd1 vssd1 vccd1 vccd1 _7940_/X sky130_fd_sc_hd__and3_1
XFILLER_48_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7871_ _7872_/B _7875_/A _7872_/A vssd1 vssd1 vccd1 vccd1 _8138_/A sky130_fd_sc_hd__o21ai_2
XFILLER_35_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6822_ _6823_/A _6823_/B vssd1 vssd1 vccd1 vccd1 _6891_/B sky130_fd_sc_hd__xnor2_1
XFILLER_90_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6753_ _6760_/A vssd1 vssd1 vccd1 vccd1 _6757_/A sky130_fd_sc_hd__inv_2
X_5704_ _5704_/A _5704_/B vssd1 vssd1 vccd1 vccd1 _6381_/B sky130_fd_sc_hd__xor2_1
XFILLER_10_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6684_ _6897_/A vssd1 vssd1 vccd1 vccd1 _7416_/A sky130_fd_sc_hd__buf_2
X_8423_ _8423_/A _8492_/B vssd1 vssd1 vccd1 vccd1 _8424_/B sky130_fd_sc_hd__xnor2_1
X_5635_ _5634_/A _5634_/C _5634_/B vssd1 vssd1 vccd1 vccd1 _5819_/D sky130_fd_sc_hd__a21oi_2
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8354_ _8354_/A _8355_/A vssd1 vssd1 vccd1 vccd1 _8358_/B sky130_fd_sc_hd__or2_1
X_5566_ _5566_/A vssd1 vssd1 vccd1 vccd1 _5680_/A sky130_fd_sc_hd__clkbuf_4
X_8285_ _8285_/A _8346_/B vssd1 vssd1 vccd1 vccd1 _8286_/B sky130_fd_sc_hd__xnor2_2
X_5497_ _8708_/Q _8666_/Q vssd1 vssd1 vccd1 vccd1 _5526_/B sky130_fd_sc_hd__xnor2_4
X_7305_ _7305_/A _7305_/B vssd1 vssd1 vccd1 vccd1 _7397_/A sky130_fd_sc_hd__xnor2_1
X_4517_ _7684_/B vssd1 vssd1 vccd1 vccd1 _4902_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_4448_ _4450_/A vssd1 vssd1 vccd1 vccd1 _4448_/Y sky130_fd_sc_hd__inv_2
X_7236_ _7236_/A _7323_/A vssd1 vssd1 vccd1 vccd1 _7237_/B sky130_fd_sc_hd__xnor2_1
XFILLER_98_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4379_ _4382_/A vssd1 vssd1 vccd1 vccd1 _4379_/Y sky130_fd_sc_hd__inv_2
X_7167_ _7167_/A _7025_/A vssd1 vssd1 vccd1 vccd1 _7219_/A sky130_fd_sc_hd__or2b_1
X_6118_ _6119_/A _6119_/B _6119_/C vssd1 vssd1 vccd1 vccd1 _6120_/A sky130_fd_sc_hd__o21a_1
XFILLER_100_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7098_ _7098_/A _7098_/B vssd1 vssd1 vccd1 vccd1 _7117_/B sky130_fd_sc_hd__xnor2_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6049_ _6049_/A vssd1 vssd1 vccd1 vccd1 _6363_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_73_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5420_ _6415_/A _6415_/B vssd1 vssd1 vccd1 vccd1 _6423_/A sky130_fd_sc_hd__and2_1
X_5351_ _8685_/Q _8684_/Q vssd1 vssd1 vccd1 vccd1 _5352_/C sky130_fd_sc_hd__nand2_1
XFILLER_99_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8070_ _8182_/B _8070_/B vssd1 vssd1 vccd1 vccd1 _8151_/B sky130_fd_sc_hd__xnor2_1
X_5282_ _5291_/B _5285_/C _5280_/X _5281_/X _5173_/B vssd1 vssd1 vccd1 vccd1 _5282_/X
+ sky130_fd_sc_hd__o32a_1
X_7021_ _7417_/A _7021_/B vssd1 vssd1 vccd1 vccd1 _7198_/C sky130_fd_sc_hd__xnor2_1
XFILLER_68_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8972_ _8972_/A _4466_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[21] sky130_fd_sc_hd__ebufn_8
X_7923_ _7998_/A _8010_/A vssd1 vssd1 vccd1 vccd1 _7928_/A sky130_fd_sc_hd__nor2_1
XFILLER_55_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7854_ _7854_/A _7854_/B vssd1 vssd1 vccd1 vccd1 _7855_/B sky130_fd_sc_hd__xor2_1
XFILLER_36_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7785_ _7719_/A _7719_/B _7784_/Y _7710_/X vssd1 vssd1 vccd1 vccd1 _7891_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_23_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6805_ _6888_/A _6805_/B vssd1 vssd1 vccd1 vccd1 _6807_/B sky130_fd_sc_hd__nor2_1
XFILLER_23_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6736_ _7685_/A _8751_/Q vssd1 vssd1 vccd1 vccd1 _6736_/X sky130_fd_sc_hd__or2b_1
X_4997_ _5225_/B _5234_/A _4980_/X _4996_/X _5130_/A vssd1 vssd1 vccd1 vccd1 _4997_/X
+ sky130_fd_sc_hd__o311a_1
X_6667_ _6694_/A _7302_/A vssd1 vssd1 vccd1 vccd1 _6799_/A sky130_fd_sc_hd__nor2_2
X_8406_ _8481_/A _8481_/B vssd1 vssd1 vccd1 vccd1 _8479_/A sky130_fd_sc_hd__nand2_1
X_5618_ _6433_/A _6653_/B vssd1 vssd1 vccd1 vccd1 _5619_/B sky130_fd_sc_hd__nor2_1
X_6598_ _6597_/A _6602_/A _6602_/B _6597_/D vssd1 vssd1 vccd1 vccd1 _6598_/X sky130_fd_sc_hd__a22o_1
X_8337_ _8337_/A _8337_/B vssd1 vssd1 vccd1 vccd1 _8338_/B sky130_fd_sc_hd__xnor2_1
X_5549_ _5917_/A _5682_/B _5853_/A _6169_/A vssd1 vssd1 vccd1 vccd1 _5549_/X sky130_fd_sc_hd__o22a_1
XFILLER_3_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8268_ _8268_/A _8268_/B _8268_/C vssd1 vssd1 vccd1 vccd1 _8280_/A sky130_fd_sc_hd__nand3_1
XFILLER_2_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8199_ _8237_/A _8238_/A vssd1 vssd1 vccd1 vccd1 _8201_/B sky130_fd_sc_hd__xnor2_1
X_8805__22 vssd1 vssd1 vccd1 vccd1 _8805__22/HI _8900_/A sky130_fd_sc_hd__conb_1
X_7219_ _7219_/A _7219_/B _7219_/C vssd1 vssd1 vccd1 vccd1 _7220_/B sky130_fd_sc_hd__and3_1
XFILLER_86_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_6_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_6_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_49_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4920_ _4920_/A _5098_/B vssd1 vssd1 vccd1 vccd1 _4956_/A sky130_fd_sc_hd__or2_1
XFILLER_33_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4851_ _4851_/A _5107_/A vssd1 vssd1 vccd1 vccd1 _4910_/B sky130_fd_sc_hd__nor2_2
X_4782_ _4549_/A _4850_/A _4779_/X _7621_/A vssd1 vssd1 vccd1 vccd1 _8664_/D sky130_fd_sc_hd__o211a_1
X_7570_ _8762_/Q _5360_/X _6569_/A _7569_/Y vssd1 vssd1 vccd1 vccd1 _8762_/D sky130_fd_sc_hd__a22o_1
X_6521_ _6521_/A _6521_/B vssd1 vssd1 vccd1 vccd1 _8743_/D sky130_fd_sc_hd__nor2_1
X_6452_ _6452_/A _6497_/B vssd1 vssd1 vccd1 vccd1 _6454_/C sky130_fd_sc_hd__nand2_1
X_5403_ _5404_/B _5403_/B vssd1 vssd1 vccd1 vccd1 _8700_/D sky130_fd_sc_hd__nor2_1
X_8122_ _8190_/A vssd1 vssd1 vccd1 vccd1 _8122_/Y sky130_fd_sc_hd__inv_2
X_6383_ _6390_/B _6383_/B _5709_/Y vssd1 vssd1 vccd1 vccd1 _6383_/X sky130_fd_sc_hd__or3b_2
X_5334_ _8683_/Q _5334_/B vssd1 vssd1 vccd1 vccd1 _5334_/X sky130_fd_sc_hd__or2_1
X_8053_ _8053_/A _8053_/B _8053_/C vssd1 vssd1 vccd1 vccd1 _8556_/A sky130_fd_sc_hd__nand3_2
X_5265_ _5291_/A _5265_/B _5265_/C _5277_/D vssd1 vssd1 vccd1 vccd1 _5265_/X sky130_fd_sc_hd__or4_1
X_7004_ _7198_/B _7004_/B vssd1 vssd1 vccd1 vccd1 _7005_/B sky130_fd_sc_hd__nand2_1
X_5196_ _4819_/X _4974_/X _5144_/X _5152_/X _5195_/X vssd1 vssd1 vccd1 vccd1 _5196_/X
+ sky130_fd_sc_hd__o41a_1
XFILLER_18_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8955_ _8955_/A _4436_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[4] sky130_fd_sc_hd__ebufn_8
X_7906_ _8439_/A _8073_/A _7917_/A vssd1 vssd1 vccd1 vccd1 _7908_/B sky130_fd_sc_hd__a21o_1
XFILLER_70_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8886_ _8886_/A _4363_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[5] sky130_fd_sc_hd__ebufn_8
X_7837_ _7892_/A _7892_/B vssd1 vssd1 vccd1 vccd1 _7866_/A sky130_fd_sc_hd__xnor2_1
XFILLER_24_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7768_ _7768_/A vssd1 vssd1 vccd1 vccd1 _8165_/B sky130_fd_sc_hd__clkbuf_2
X_7699_ _8772_/Q _8669_/Q vssd1 vssd1 vccd1 vccd1 _7699_/X sky130_fd_sc_hd__and2b_1
X_6719_ _6713_/A _6714_/A _6713_/B vssd1 vssd1 vccd1 vccd1 _7137_/A sky130_fd_sc_hd__a21bo_1
XFILLER_50_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5050_ _5156_/A _5077_/C _5263_/C _5050_/D vssd1 vssd1 vccd1 vccd1 _5051_/D sky130_fd_sc_hd__or4_1
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8796__13 vssd1 vssd1 vccd1 vccd1 _8796__13/HI _8891_/A sky130_fd_sc_hd__conb_1
XFILLER_38_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5952_ _5953_/A _5953_/B vssd1 vssd1 vccd1 vccd1 _6047_/A sky130_fd_sc_hd__nor2_1
XFILLER_80_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8740_ _8742_/CLK _8740_/D vssd1 vssd1 vccd1 vccd1 _8740_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4903_ _5082_/B _4912_/B vssd1 vssd1 vccd1 vccd1 _5119_/A sky130_fd_sc_hd__nor2_2
X_5883_ _5883_/A _5881_/B vssd1 vssd1 vccd1 vccd1 _6128_/A sky130_fd_sc_hd__or2b_1
X_8671_ _8771_/CLK _8671_/D vssd1 vssd1 vccd1 vccd1 _8671_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_33_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7622_ _7622_/A _7622_/B vssd1 vssd1 vccd1 vccd1 _7649_/B sky130_fd_sc_hd__nor2_2
X_4834_ _5184_/B vssd1 vssd1 vccd1 vccd1 _5148_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_21_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4765_ _5100_/A _4767_/B vssd1 vssd1 vccd1 vccd1 _4765_/X sky130_fd_sc_hd__and2_1
X_7553_ _7541_/X _7552_/X _5491_/X _8758_/Q vssd1 vssd1 vccd1 vccd1 _8758_/D sky130_fd_sc_hd__o2bb2a_1
X_6504_ _6506_/B _6506_/C _6465_/X vssd1 vssd1 vccd1 vccd1 _6504_/Y sky130_fd_sc_hd__o21ai_1
X_7484_ _7482_/X _7483_/X _7484_/S vssd1 vssd1 vccd1 vccd1 _7486_/A sky130_fd_sc_hd__mux2_1
X_4696_ _4720_/A vssd1 vssd1 vccd1 vccd1 _4697_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6435_ _7589_/A _6435_/B _6435_/C vssd1 vssd1 vccd1 vccd1 _6436_/A sky130_fd_sc_hd__and3_1
X_6366_ _6365_/B _6365_/C _6365_/A vssd1 vssd1 vccd1 vccd1 _6366_/Y sky130_fd_sc_hd__o21ai_1
X_8105_ _8568_/A _8497_/A vssd1 vssd1 vccd1 vccd1 _8343_/A sky130_fd_sc_hd__or2_2
X_5317_ _8717_/Q _5307_/X _5316_/X _5311_/X vssd1 vssd1 vccd1 vccd1 _8675_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6297_ _6297_/A _6361_/A vssd1 vssd1 vccd1 vccd1 _6360_/A sky130_fd_sc_hd__nand2_1
XFILLER_102_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8036_ _8036_/A _8036_/B vssd1 vssd1 vccd1 vccd1 _8036_/Y sky130_fd_sc_hd__nand2_1
XFILLER_102_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5248_ _5133_/Y _5245_/Y _5246_/Y _5247_/X vssd1 vssd1 vccd1 vccd1 _5248_/X sky130_fd_sc_hd__a211o_1
XFILLER_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5179_ _5281_/A _5179_/B _5179_/C _5179_/D vssd1 vssd1 vccd1 vccd1 _5179_/X sky130_fd_sc_hd__or4_1
XFILLER_56_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8938_ _8938_/A _4427_/Y vssd1 vssd1 vccd1 vccd1 io_out[25] sky130_fd_sc_hd__ebufn_8
XFILLER_83_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8880__97 vssd1 vssd1 vccd1 vccd1 _8880__97/HI _8704_/D sky130_fd_sc_hd__conb_1
XFILLER_86_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4550_ _4550_/A vssd1 vssd1 vccd1 vccd1 _8925_/A sky130_fd_sc_hd__clkbuf_1
X_4481_ _4481_/A vssd1 vssd1 vccd1 vccd1 _4486_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6220_ _6162_/A _6162_/B _6219_/X vssd1 vssd1 vccd1 vccd1 _6288_/A sky130_fd_sc_hd__a21oi_1
X_6151_ _6224_/A _6224_/B vssd1 vssd1 vccd1 vccd1 _6152_/B sky130_fd_sc_hd__xor2_1
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5102_ _5098_/X _5099_/X _5221_/A _5215_/B _5188_/D vssd1 vssd1 vccd1 vccd1 _5102_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6082_ _5995_/A _5995_/B _6081_/X vssd1 vssd1 vccd1 vccd1 _6087_/A sky130_fd_sc_hd__a21oi_2
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5033_ _5033_/A _5033_/B vssd1 vssd1 vccd1 vccd1 _5228_/B sky130_fd_sc_hd__or2_2
XFILLER_65_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6984_ _6984_/A _6983_/A vssd1 vssd1 vccd1 vccd1 _6984_/X sky130_fd_sc_hd__or2b_1
X_5935_ _6011_/A _6011_/B vssd1 vssd1 vccd1 vccd1 _5939_/A sky130_fd_sc_hd__xnor2_1
X_8723_ _8723_/CLK _8723_/D vssd1 vssd1 vccd1 vccd1 _8723_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5866_ _5942_/A _5866_/B vssd1 vssd1 vccd1 vccd1 _5867_/C sky130_fd_sc_hd__xor2_1
XFILLER_80_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8654_ _8778_/CLK _8654_/D vssd1 vssd1 vccd1 vccd1 _8654_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4817_ _4817_/A vssd1 vssd1 vccd1 vccd1 _8671_/D sky130_fd_sc_hd__clkbuf_1
X_7605_ _7602_/A _7622_/B _8621_/B vssd1 vssd1 vccd1 vccd1 _7606_/C sky130_fd_sc_hd__a21bo_1
XFILLER_21_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5797_ _5766_/A _5921_/B _5666_/B _5796_/X vssd1 vssd1 vccd1 vccd1 _5799_/B sky130_fd_sc_hd__a31oi_1
X_8585_ _7624_/X _8573_/X _8583_/X _8584_/Y vssd1 vssd1 vccd1 vccd1 _8777_/D sky130_fd_sc_hd__a31oi_1
X_4748_ _4748_/A vssd1 vssd1 vccd1 vccd1 _8658_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7536_ _7536_/A _7536_/B vssd1 vssd1 vccd1 vccd1 _7537_/B sky130_fd_sc_hd__and2_1
X_4679_ _4679_/A _4679_/B _4679_/C vssd1 vssd1 vccd1 vccd1 _4680_/A sky130_fd_sc_hd__and3_1
X_7467_ _7467_/A _7467_/B vssd1 vssd1 vccd1 vccd1 _7470_/A sky130_fd_sc_hd__or2_1
X_6418_ _5421_/Y _6423_/B _6417_/Y _5443_/B vssd1 vssd1 vccd1 vccd1 _6418_/X sky130_fd_sc_hd__a211o_1
X_7398_ _7316_/A _7316_/B _7397_/X vssd1 vssd1 vccd1 vccd1 _7399_/B sky130_fd_sc_hd__a21oi_2
X_6349_ _6349_/A _6349_/B vssd1 vssd1 vccd1 vccd1 _6354_/A sky130_fd_sc_hd__xnor2_1
XFILLER_88_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8019_ _8059_/A _8018_/C _8018_/A vssd1 vssd1 vccd1 vccd1 _8020_/C sky130_fd_sc_hd__a21o_1
XFILLER_91_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5720_ _5986_/A _5720_/B vssd1 vssd1 vccd1 vccd1 _5720_/Y sky130_fd_sc_hd__nand2_1
X_5651_ _5544_/A _5541_/Y _5544_/B _5542_/A vssd1 vssd1 vccd1 vccd1 _5652_/B sky130_fd_sc_hd__a31o_1
X_8370_ _8370_/A _8370_/B vssd1 vssd1 vccd1 vccd1 _8371_/B sky130_fd_sc_hd__nor2_1
X_5582_ _5701_/B vssd1 vssd1 vccd1 vccd1 _6004_/A sky130_fd_sc_hd__clkbuf_2
X_4602_ _6563_/B vssd1 vssd1 vccd1 vccd1 _4807_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7321_ _7321_/A _7321_/B vssd1 vssd1 vccd1 vccd1 _7322_/B sky130_fd_sc_hd__xnor2_2
X_4533_ _8662_/Q vssd1 vssd1 vccd1 vccd1 _4878_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_7252_ _7346_/A _7252_/B vssd1 vssd1 vccd1 vccd1 _7348_/B sky130_fd_sc_hd__nand2_1
XFILLER_89_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6203_ _6278_/A _6203_/B _6278_/B vssd1 vssd1 vccd1 vccd1 _6204_/B sky130_fd_sc_hd__and3_1
X_4464_ _4468_/A vssd1 vssd1 vccd1 vccd1 _4464_/Y sky130_fd_sc_hd__inv_2
X_4395_ _4395_/A vssd1 vssd1 vccd1 vccd1 _4400_/A sky130_fd_sc_hd__buf_6
X_7183_ _7285_/B _7183_/B vssd1 vssd1 vccd1 vccd1 _7288_/B sky130_fd_sc_hd__or2_1
X_6134_ _6134_/A _6134_/B vssd1 vssd1 vccd1 vccd1 _6134_/Y sky130_fd_sc_hd__nor2_1
XFILLER_58_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6065_ _6065_/A _6065_/B vssd1 vssd1 vccd1 vccd1 _6104_/A sky130_fd_sc_hd__xor2_2
XFILLER_58_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5016_ _5155_/C _5285_/B vssd1 vssd1 vccd1 vccd1 _5174_/B sky130_fd_sc_hd__or2_2
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6967_ _6967_/A _6967_/B vssd1 vssd1 vccd1 vccd1 _6967_/X sky130_fd_sc_hd__xor2_1
X_5918_ _6059_/A _6230_/A vssd1 vssd1 vccd1 vccd1 _5918_/X sky130_fd_sc_hd__and2_1
X_8706_ _8720_/CLK _8706_/D vssd1 vssd1 vccd1 vccd1 _8706_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6898_ _6898_/A _7036_/A vssd1 vssd1 vccd1 vccd1 _7282_/A sky130_fd_sc_hd__or2_2
X_5849_ _5779_/A _5849_/B vssd1 vssd1 vccd1 vccd1 _5936_/A sky130_fd_sc_hd__and2b_1
XFILLER_21_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8637_ _8732_/CLK _8637_/D vssd1 vssd1 vccd1 vccd1 _8637_/Q sky130_fd_sc_hd__dfxtp_1
X_8568_ _8568_/A _8568_/B _8568_/C _8568_/D vssd1 vssd1 vccd1 vccd1 _8568_/X sky130_fd_sc_hd__and4_1
XFILLER_5_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7519_ _7519_/A _7519_/B vssd1 vssd1 vccd1 vccd1 _7539_/A sky130_fd_sc_hd__xnor2_1
X_8499_ _8499_/A _8499_/B vssd1 vssd1 vccd1 vccd1 _8500_/B sky130_fd_sc_hd__xnor2_1
X_8850__67 vssd1 vssd1 vccd1 vccd1 _8850__67/HI _8959_/A sky130_fd_sc_hd__conb_1
XFILLER_57_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7870_ _7891_/A _7891_/B vssd1 vssd1 vccd1 vccd1 _7872_/A sky130_fd_sc_hd__xor2_1
XFILLER_63_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6821_ _6953_/A _6821_/B vssd1 vssd1 vccd1 vccd1 _6823_/B sky130_fd_sc_hd__nor2_1
XFILLER_35_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6752_ _6752_/A _6752_/B vssd1 vssd1 vccd1 vccd1 _6760_/A sky130_fd_sc_hd__nor2_1
X_5703_ _6378_/C _6070_/A vssd1 vssd1 vccd1 vccd1 _6377_/B sky130_fd_sc_hd__nor2_1
X_6683_ _7363_/B _7379_/B vssd1 vssd1 vccd1 vccd1 _6897_/A sky130_fd_sc_hd__or2_1
X_8422_ _8422_/A _8422_/B vssd1 vssd1 vccd1 vccd1 _8492_/B sky130_fd_sc_hd__xor2_1
X_5634_ _5634_/A _5634_/B _5634_/C vssd1 vssd1 vccd1 vccd1 _5819_/C sky130_fd_sc_hd__and3_1
X_8353_ _8327_/A _8418_/A _8352_/Y _8336_/A vssd1 vssd1 vccd1 vccd1 _8353_/X sky130_fd_sc_hd__o22a_1
X_5565_ _8655_/Q _8718_/Q vssd1 vssd1 vccd1 vccd1 _5566_/A sky130_fd_sc_hd__or2b_1
X_7304_ _7382_/A _7304_/B vssd1 vssd1 vccd1 vccd1 _7305_/B sky130_fd_sc_hd__xnor2_1
X_8284_ _8284_/A _8284_/B vssd1 vssd1 vccd1 vccd1 _8346_/B sky130_fd_sc_hd__xor2_1
X_5496_ _5773_/A vssd1 vssd1 vccd1 vccd1 _6378_/A sky130_fd_sc_hd__clkbuf_2
X_4516_ _8668_/Q vssd1 vssd1 vccd1 vccd1 _7684_/B sky130_fd_sc_hd__buf_2
X_4447_ _4450_/A vssd1 vssd1 vccd1 vccd1 _4447_/Y sky130_fd_sc_hd__clkinv_4
X_7235_ _7235_/A _7235_/B vssd1 vssd1 vccd1 vccd1 _7323_/A sky130_fd_sc_hd__xnor2_1
XFILLER_104_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7166_ _7061_/A _7061_/B _7165_/Y vssd1 vssd1 vccd1 vccd1 _7241_/A sky130_fd_sc_hd__a21bo_1
X_6117_ _6162_/A _6117_/B vssd1 vssd1 vccd1 vccd1 _6119_/C sky130_fd_sc_hd__and2b_1
X_4378_ _4382_/A vssd1 vssd1 vccd1 vccd1 _4378_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7097_ _7097_/A _7097_/B vssd1 vssd1 vccd1 vccd1 _7157_/A sky130_fd_sc_hd__xor2_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6048_ _6129_/A _6129_/B vssd1 vssd1 vccd1 vccd1 _6049_/A sky130_fd_sc_hd__and2_1
XFILLER_54_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7999_ _7999_/A vssd1 vssd1 vccd1 vccd1 _7999_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_81_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_8_0_wb_clk_i clkbuf_4_9_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _8763_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5350_ _5355_/A vssd1 vssd1 vccd1 vccd1 _5409_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_99_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5281_ _5281_/A _5281_/B _5285_/B vssd1 vssd1 vccd1 vccd1 _5281_/X sky130_fd_sc_hd__or3_1
XFILLER_4_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7020_ _7020_/A _7020_/B vssd1 vssd1 vccd1 vccd1 _7021_/B sky130_fd_sc_hd__nand2_2
XFILLER_101_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8971_ _8971_/A _4465_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[20] sky130_fd_sc_hd__ebufn_8
XFILLER_67_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7922_ _7921_/B _7921_/C _7921_/A vssd1 vssd1 vccd1 vccd1 _7930_/B sky130_fd_sc_hd__a21o_1
XFILLER_36_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7853_ _7959_/A _7959_/B vssd1 vssd1 vccd1 vccd1 _7860_/A sky130_fd_sc_hd__xor2_1
XFILLER_63_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7784_ _7784_/A _7784_/B vssd1 vssd1 vccd1 vccd1 _7784_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6804_ _6804_/A _6804_/B vssd1 vssd1 vccd1 vccd1 _6805_/B sky130_fd_sc_hd__and2_1
X_4996_ _4990_/X _4995_/X _4819_/X vssd1 vssd1 vccd1 vccd1 _4996_/X sky130_fd_sc_hd__a21o_1
XFILLER_51_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6735_ _6735_/A _6735_/B vssd1 vssd1 vccd1 vccd1 _6764_/B sky130_fd_sc_hd__nor2_4
X_6666_ _7034_/A vssd1 vssd1 vccd1 vccd1 _7302_/A sky130_fd_sc_hd__clkbuf_2
X_8405_ _8405_/A _8408_/B vssd1 vssd1 vccd1 vccd1 _8481_/B sky130_fd_sc_hd__xnor2_2
X_5617_ _5617_/A _6653_/B vssd1 vssd1 vccd1 vccd1 _5619_/A sky130_fd_sc_hd__and2_1
X_6597_ _6597_/A _6602_/A _6602_/B _6597_/D vssd1 vssd1 vccd1 vccd1 _6599_/A sky130_fd_sc_hd__and4_1
X_8336_ _8336_/A _8352_/A vssd1 vssd1 vccd1 vccd1 _8337_/B sky130_fd_sc_hd__xnor2_1
X_5548_ _5917_/A _6169_/A vssd1 vssd1 vccd1 vccd1 _5662_/B sky130_fd_sc_hd__nor2_1
X_8267_ _8386_/B _8266_/C _8266_/A vssd1 vssd1 vccd1 vccd1 _8268_/C sky130_fd_sc_hd__a21o_1
XFILLER_78_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7218_ _7219_/A _7219_/B _7219_/C vssd1 vssd1 vccd1 vccd1 _7220_/A sky130_fd_sc_hd__a21oi_1
X_5479_ _5480_/A _5485_/S _5480_/C _5484_/B vssd1 vssd1 vccd1 vccd1 _5481_/A sky130_fd_sc_hd__a22o_1
X_8198_ _8198_/A _8343_/A _8420_/A vssd1 vssd1 vccd1 vccd1 _8238_/A sky130_fd_sc_hd__and3_1
X_7149_ _7536_/A _7536_/B vssd1 vssd1 vccd1 vccd1 _7537_/A sky130_fd_sc_hd__nor2_1
XFILLER_100_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8820__37 vssd1 vssd1 vccd1 vccd1 _8820__37/HI _8915_/A sky130_fd_sc_hd__conb_1
XFILLER_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4850_ _4850_/A _4901_/B _4850_/C vssd1 vssd1 vccd1 vccd1 _5107_/A sky130_fd_sc_hd__and3_1
XFILLER_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4781_ _5335_/A vssd1 vssd1 vccd1 vccd1 _7621_/A sky130_fd_sc_hd__clkbuf_4
X_6520_ _8743_/Q _6519_/B _6483_/X vssd1 vssd1 vccd1 vccd1 _6521_/B sky130_fd_sc_hd__o21ai_1
X_6451_ _8735_/Q vssd1 vssd1 vccd1 vccd1 _6497_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6382_ _5710_/A _6389_/B _5807_/X vssd1 vssd1 vccd1 vccd1 _6383_/B sky130_fd_sc_hd__a21bo_1
X_5402_ _8700_/Q _5400_/A _5392_/X vssd1 vssd1 vccd1 vccd1 _5403_/B sky130_fd_sc_hd__o21ai_1
X_8121_ _8289_/B _8121_/B vssd1 vssd1 vccd1 vccd1 _8124_/A sky130_fd_sc_hd__or2_1
X_5333_ _8757_/Q _5320_/A _5332_/X _5324_/X vssd1 vssd1 vccd1 vccd1 _8682_/D sky130_fd_sc_hd__o211a_1
XFILLER_102_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8052_ _8055_/A _8051_/C _8051_/A vssd1 vssd1 vccd1 vccd1 _8053_/C sky130_fd_sc_hd__o21ai_1
X_5264_ _5264_/A _5283_/B vssd1 vssd1 vccd1 vccd1 _5277_/D sky130_fd_sc_hd__or2_1
XFILLER_87_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7003_ _7380_/A _7004_/B vssd1 vssd1 vccd1 vccd1 _7288_/A sky130_fd_sc_hd__or2_2
X_5195_ _5170_/X _5181_/Y _5194_/X _5130_/A vssd1 vssd1 vccd1 vccd1 _5195_/X sky130_fd_sc_hd__a31o_1
XFILLER_68_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8954_ _8954_/A _4437_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[3] sky130_fd_sc_hd__ebufn_8
XFILLER_83_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7905_ _8273_/A _8172_/A vssd1 vssd1 vccd1 vccd1 _7917_/A sky130_fd_sc_hd__nor2_2
X_8885_ _8885_/A _4362_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[4] sky130_fd_sc_hd__ebufn_8
XFILLER_36_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7836_ _8261_/A _8568_/D _7836_/C vssd1 vssd1 vccd1 vccd1 _7892_/B sky130_fd_sc_hd__or3_1
XFILLER_24_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7767_ _7913_/A _7902_/A vssd1 vssd1 vccd1 vccd1 _7880_/A sky130_fd_sc_hd__nor2_1
X_4979_ _5078_/B _5149_/B vssd1 vssd1 vccd1 vccd1 _5096_/B sky130_fd_sc_hd__or2_2
X_7698_ _7688_/A _7688_/B _7686_/B _7684_/X vssd1 vssd1 vccd1 vccd1 _7702_/A sky130_fd_sc_hd__a31o_1
X_6718_ _7392_/A _6957_/A vssd1 vssd1 vccd1 vccd1 _6721_/A sky130_fd_sc_hd__xnor2_1
X_6649_ _6694_/A _6810_/A vssd1 vssd1 vccd1 vccd1 _6924_/A sky130_fd_sc_hd__or2_2
X_8319_ _8303_/B _8305_/B _8303_/A vssd1 vssd1 vccd1 vccd1 _8405_/A sky130_fd_sc_hd__o21ba_1
XFILLER_3_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5951_ _6044_/A _5951_/B vssd1 vssd1 vccd1 vccd1 _5953_/B sky130_fd_sc_hd__nand2_1
XFILLER_52_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4902_ _4874_/B _4902_/B _4902_/C vssd1 vssd1 vccd1 vccd1 _5009_/C sky130_fd_sc_hd__and3b_2
X_8670_ _8758_/CLK _8670_/D vssd1 vssd1 vccd1 vccd1 _8670_/Q sky130_fd_sc_hd__dfxtp_1
X_5882_ _5961_/B vssd1 vssd1 vccd1 vccd1 _6370_/A sky130_fd_sc_hd__buf_2
X_7621_ _7621_/A _7621_/B vssd1 vssd1 vccd1 vccd1 _8767_/D sky130_fd_sc_hd__nand2_1
XFILLER_60_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4833_ _5206_/A vssd1 vssd1 vccd1 vccd1 _5184_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_7552_ _7552_/A _7552_/B _7552_/C vssd1 vssd1 vccd1 vccd1 _7552_/X sky130_fd_sc_hd__or3_1
X_4764_ _4702_/A _4702_/B _4818_/B _5259_/D vssd1 vssd1 vccd1 vccd1 _4767_/B sky130_fd_sc_hd__and4bb_2
X_7483_ _7482_/B _7483_/B vssd1 vssd1 vccd1 vccd1 _7483_/X sky130_fd_sc_hd__and2b_1
X_6503_ _6506_/C _6503_/B vssd1 vssd1 vccd1 vccd1 _8737_/D sky130_fd_sc_hd__nor2_1
X_4695_ _5181_/A _4695_/B vssd1 vssd1 vccd1 vccd1 _4702_/B sky130_fd_sc_hd__nand2_1
X_6434_ _5462_/X _6432_/X _8724_/Q vssd1 vssd1 vccd1 vccd1 _6435_/C sky130_fd_sc_hd__a21o_1
X_6365_ _6365_/A _6365_/B _6365_/C vssd1 vssd1 vccd1 vccd1 _6365_/X sky130_fd_sc_hd__or3_1
X_6296_ _6296_/A _6296_/B vssd1 vssd1 vccd1 vccd1 _6361_/A sky130_fd_sc_hd__or2_1
X_8104_ _8348_/B vssd1 vssd1 vccd1 vccd1 _8497_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5316_ _8675_/Q _5326_/B vssd1 vssd1 vccd1 vccd1 _5316_/X sky130_fd_sc_hd__or2_1
XFILLER_88_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8035_ _8114_/A _8114_/B vssd1 vssd1 vccd1 vccd1 _8119_/A sky130_fd_sc_hd__xnor2_1
X_5247_ _5300_/B _5247_/B vssd1 vssd1 vccd1 vccd1 _5247_/X sky130_fd_sc_hd__and2_1
XFILLER_0_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5178_ _5192_/A _5178_/B vssd1 vssd1 vccd1 vccd1 _5179_/D sky130_fd_sc_hd__or2_1
X_8937_ _8937_/A _4425_/Y vssd1 vssd1 vccd1 vccd1 io_out[24] sky130_fd_sc_hd__ebufn_8
XFILLER_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7819_ _7819_/A _7819_/B vssd1 vssd1 vccd1 vccd1 _7895_/C sky130_fd_sc_hd__xor2_1
XFILLER_12_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4480_ _4480_/A vssd1 vssd1 vccd1 vccd1 _4480_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8856__73 vssd1 vssd1 vccd1 vccd1 _8856__73/HI _8965_/A sky130_fd_sc_hd__conb_1
X_6150_ _5928_/B _6150_/B _6227_/B vssd1 vssd1 vccd1 vccd1 _6224_/B sky130_fd_sc_hd__and3b_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5101_ _5221_/B _5101_/B vssd1 vssd1 vccd1 vccd1 _5188_/D sky130_fd_sc_hd__or2_2
X_6081_ _6081_/A _6193_/A _6274_/B vssd1 vssd1 vccd1 vccd1 _6081_/X sky130_fd_sc_hd__and3_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_10_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8758_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_97_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5032_ _5040_/B _5032_/B vssd1 vssd1 vccd1 vccd1 _5036_/A sky130_fd_sc_hd__nor2_1
XFILLER_38_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6983_ _6983_/A _6984_/A vssd1 vssd1 vccd1 vccd1 _7090_/B sky130_fd_sc_hd__xnor2_1
XFILLER_25_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5934_ _5934_/A _5934_/B vssd1 vssd1 vccd1 vccd1 _6011_/B sky130_fd_sc_hd__nor2_1
X_8722_ _8723_/CLK _8722_/D vssd1 vssd1 vccd1 vccd1 _8722_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5865_ _5786_/A _5786_/B _5864_/Y vssd1 vssd1 vccd1 vccd1 _5866_/B sky130_fd_sc_hd__o21ai_1
XFILLER_80_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8653_ _8778_/CLK _8653_/D vssd1 vssd1 vccd1 vccd1 _8653_/Q sky130_fd_sc_hd__dfxtp_1
X_7604_ _7599_/X _7602_/X _8784_/Q _8626_/A vssd1 vssd1 vccd1 vccd1 _7606_/B sky130_fd_sc_hd__a211o_1
X_4816_ _5335_/A _4816_/B vssd1 vssd1 vccd1 vccd1 _4817_/A sky130_fd_sc_hd__and2_1
X_5796_ _5764_/A _5796_/B vssd1 vssd1 vccd1 vccd1 _5796_/X sky130_fd_sc_hd__and2b_1
X_8584_ _8588_/A _8777_/Q vssd1 vssd1 vccd1 vccd1 _8584_/Y sky130_fd_sc_hd__nor2_1
X_4747_ _4751_/B _4747_/B _4747_/C vssd1 vssd1 vccd1 vccd1 _4748_/A sky130_fd_sc_hd__and3b_1
X_7535_ _7535_/A _7552_/A _7552_/B vssd1 vssd1 vccd1 vccd1 _7535_/X sky130_fd_sc_hd__or3_1
X_4678_ _8650_/Q _4678_/B vssd1 vssd1 vccd1 vccd1 _4679_/C sky130_fd_sc_hd__nand2_1
X_7466_ _7465_/A _7465_/B _7465_/C vssd1 vssd1 vccd1 vccd1 _7467_/B sky130_fd_sc_hd__a21oi_1
X_7397_ _7397_/A _7397_/B vssd1 vssd1 vccd1 vccd1 _7397_/X sky130_fd_sc_hd__and2_1
X_6417_ _5421_/Y _6416_/B _6416_/A vssd1 vssd1 vccd1 vccd1 _6417_/Y sky130_fd_sc_hd__a21oi_1
X_6348_ _6348_/A _6348_/B vssd1 vssd1 vccd1 vccd1 _6349_/B sky130_fd_sc_hd__xnor2_1
XFILLER_88_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6279_ _6279_/A _6279_/B vssd1 vssd1 vccd1 vccd1 _6280_/B sky130_fd_sc_hd__nor2_1
XFILLER_88_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8018_ _8018_/A _8059_/A _8018_/C vssd1 vssd1 vccd1 vccd1 _8059_/B sky130_fd_sc_hd__nand3_1
XFILLER_29_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8786__3 vssd1 vssd1 vccd1 vccd1 _8786__3/HI _8881_/A sky130_fd_sc_hd__conb_1
XFILLER_21_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5650_ _5925_/A _5650_/B vssd1 vssd1 vccd1 vccd1 _5769_/A sky130_fd_sc_hd__nand2_1
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4601_ input2/X vssd1 vssd1 vccd1 vccd1 _6563_/B sky130_fd_sc_hd__buf_2
X_5581_ _5680_/A _5680_/B vssd1 vssd1 vccd1 vccd1 _5701_/B sky130_fd_sc_hd__xor2_4
X_7320_ _7320_/A _7320_/B vssd1 vssd1 vccd1 vccd1 _7321_/B sky130_fd_sc_hd__xnor2_2
XFILLER_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4532_ _4774_/A vssd1 vssd1 vccd1 vccd1 _4872_/B sky130_fd_sc_hd__clkbuf_1
X_4463_ _4481_/A vssd1 vssd1 vccd1 vccd1 _4468_/A sky130_fd_sc_hd__buf_2
X_7251_ _7251_/A _7243_/A vssd1 vssd1 vccd1 vccd1 _7348_/A sky130_fd_sc_hd__or2b_1
XFILLER_104_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6202_ _6278_/A _6203_/B _6278_/B vssd1 vssd1 vccd1 vccd1 _6204_/A sky130_fd_sc_hd__a21oi_1
X_4394_ _4394_/A vssd1 vssd1 vccd1 vccd1 _4394_/Y sky130_fd_sc_hd__inv_2
X_7182_ _7182_/A _7229_/A vssd1 vssd1 vccd1 vccd1 _7183_/B sky130_fd_sc_hd__and2_1
X_6133_ _6363_/A _6365_/B _6363_/B vssd1 vssd1 vccd1 vccd1 _6360_/C sky130_fd_sc_hd__o21ai_1
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6064_ _6064_/A _6064_/B vssd1 vssd1 vccd1 vccd1 _6065_/B sky130_fd_sc_hd__xnor2_1
XFILLER_85_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5015_ _5108_/B vssd1 vssd1 vccd1 vccd1 _5285_/B sky130_fd_sc_hd__clkbuf_2
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6966_ _7141_/A _6966_/B vssd1 vssd1 vccd1 vccd1 _6968_/B sky130_fd_sc_hd__or2_1
X_5917_ _5917_/A _6165_/B vssd1 vssd1 vccd1 vccd1 _6230_/A sky130_fd_sc_hd__or2_2
X_8705_ _8720_/CLK _8705_/D vssd1 vssd1 vccd1 vccd1 _8705_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6897_ _6897_/A _7392_/A vssd1 vssd1 vccd1 vccd1 _7001_/A sky130_fd_sc_hd__or2_1
XFILLER_42_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5848_ _5887_/B _5847_/C _5847_/A vssd1 vssd1 vccd1 vccd1 _5867_/B sky130_fd_sc_hd__a21oi_1
X_8636_ _8732_/CLK _8636_/D vssd1 vssd1 vccd1 vccd1 _8636_/Q sky130_fd_sc_hd__dfxtp_1
X_5779_ _5779_/A _5849_/B vssd1 vssd1 vccd1 vccd1 _5864_/B sky130_fd_sc_hd__xnor2_1
X_8567_ _8567_/A _8567_/B vssd1 vssd1 vccd1 vccd1 _8567_/X sky130_fd_sc_hd__or2_1
XFILLER_5_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7518_ _7518_/A _7518_/B vssd1 vssd1 vccd1 vccd1 _7548_/A sky130_fd_sc_hd__nand2_1
X_8498_ _8496_/S _8357_/A _8498_/S vssd1 vssd1 vccd1 vccd1 _8499_/B sky130_fd_sc_hd__mux2_1
X_7449_ _7485_/B _7449_/B vssd1 vssd1 vccd1 vccd1 _7454_/A sky130_fd_sc_hd__xnor2_1
XFILLER_89_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8826__43 vssd1 vssd1 vccd1 vccd1 _8826__43/HI _8921_/A sky130_fd_sc_hd__conb_1
XFILLER_4_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6820_ _6820_/A _6820_/B vssd1 vssd1 vccd1 vccd1 _6821_/B sky130_fd_sc_hd__and2_1
XFILLER_23_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6751_ _6851_/A _8671_/Q vssd1 vssd1 vccd1 vccd1 _6752_/B sky130_fd_sc_hd__nor2_1
X_5702_ _5702_/A _5702_/B vssd1 vssd1 vccd1 vccd1 _6070_/A sky130_fd_sc_hd__nor2_1
Xclkbuf_1_1_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
X_6682_ _7181_/B vssd1 vssd1 vccd1 vccd1 _6682_/Y sky130_fd_sc_hd__inv_2
X_8421_ _8421_/A _8494_/B vssd1 vssd1 vccd1 vccd1 _8422_/B sky130_fd_sc_hd__xnor2_1
X_5633_ _5824_/B vssd1 vssd1 vccd1 vccd1 _6068_/B sky130_fd_sc_hd__clkbuf_2
X_8352_ _8352_/A vssd1 vssd1 vccd1 vccd1 _8352_/Y sky130_fd_sc_hd__inv_2
X_5564_ _5564_/A _5564_/B vssd1 vssd1 vccd1 vccd1 _5585_/A sky130_fd_sc_hd__nor2_2
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7303_ _7303_/A _7377_/A vssd1 vssd1 vccd1 vccd1 _7304_/B sky130_fd_sc_hd__xnor2_1
X_4515_ _7700_/A vssd1 vssd1 vccd1 vccd1 _4804_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_8283_ _8364_/A _8364_/B vssd1 vssd1 vccd1 vccd1 _8284_/B sky130_fd_sc_hd__xor2_1
X_5495_ _5552_/A _5552_/B vssd1 vssd1 vccd1 vccd1 _5773_/A sky130_fd_sc_hd__and2_2
XFILLER_104_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4446_ _4450_/A vssd1 vssd1 vccd1 vccd1 _4446_/Y sky130_fd_sc_hd__inv_2
X_7234_ _7336_/A _7336_/B vssd1 vssd1 vccd1 vccd1 _7235_/B sky130_fd_sc_hd__xnor2_1
X_4377_ _4395_/A vssd1 vssd1 vccd1 vccd1 _4382_/A sky130_fd_sc_hd__clkbuf_2
X_7165_ _7165_/A _7165_/B vssd1 vssd1 vccd1 vccd1 _7165_/Y sky130_fd_sc_hd__nand2_1
X_6116_ _6116_/A _6116_/B vssd1 vssd1 vccd1 vccd1 _6117_/B sky130_fd_sc_hd__nand2_1
XFILLER_98_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7096_ _7096_/A _7096_/B _7096_/C vssd1 vssd1 vccd1 vccd1 _7528_/B sky130_fd_sc_hd__nand3_2
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6047_ _6047_/A _6047_/B vssd1 vssd1 vccd1 vccd1 _6129_/B sky130_fd_sc_hd__xor2_1
XFILLER_73_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7998_ _7998_/A _8273_/B vssd1 vssd1 vccd1 vccd1 _7999_/A sky130_fd_sc_hd__nor2_1
XFILLER_26_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6949_ _6949_/A _6949_/B vssd1 vssd1 vccd1 vccd1 _7049_/B sky130_fd_sc_hd__or2_1
XFILLER_41_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8619_ _8619_/A _8627_/S vssd1 vssd1 vccd1 vccd1 _8623_/A sky130_fd_sc_hd__or2b_1
XFILLER_22_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5280_ _5280_/A _5285_/A _5141_/C vssd1 vssd1 vccd1 vccd1 _5280_/X sky130_fd_sc_hd__or3b_1
XFILLER_99_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8970_ _8970_/A _4464_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[19] sky130_fd_sc_hd__ebufn_8
XFILLER_67_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7921_ _7921_/A _7921_/B _7921_/C vssd1 vssd1 vccd1 vccd1 _7930_/A sky130_fd_sc_hd__nand3_1
XFILLER_82_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7852_ _8325_/A _7710_/X _7784_/Y _7711_/A vssd1 vssd1 vccd1 vccd1 _7959_/B sky130_fd_sc_hd__a211o_1
XFILLER_51_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7783_ _7783_/A _7783_/B vssd1 vssd1 vccd1 vccd1 _7784_/B sky130_fd_sc_hd__xnor2_1
XFILLER_51_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6803_ _6804_/A _6804_/B vssd1 vssd1 vccd1 vccd1 _6888_/A sky130_fd_sc_hd__nor2_2
X_4995_ _4995_/A _5007_/A _4995_/C _4995_/D vssd1 vssd1 vccd1 vccd1 _4995_/X sky130_fd_sc_hd__or4_1
X_6734_ _8751_/Q _7685_/A vssd1 vssd1 vccd1 vccd1 _6735_/B sky130_fd_sc_hd__and2b_1
XFILLER_23_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8404_ _8407_/B _8404_/B vssd1 vssd1 vccd1 vccd1 _8408_/B sky130_fd_sc_hd__xnor2_1
X_6665_ _6674_/B _6678_/A _6674_/D _7363_/A vssd1 vssd1 vccd1 vccd1 _7034_/A sky130_fd_sc_hd__a31o_2
X_5616_ _5608_/A _5608_/B _5615_/X vssd1 vssd1 vccd1 vccd1 _5620_/B sky130_fd_sc_hd__a21oi_1
X_6596_ _6758_/A _8747_/Q vssd1 vssd1 vccd1 vccd1 _6597_/D sky130_fd_sc_hd__or2_1
X_8335_ _8335_/A _8335_/B vssd1 vssd1 vccd1 vccd1 _8337_/A sky130_fd_sc_hd__xor2_1
X_5547_ _5547_/A _5547_/B vssd1 vssd1 vccd1 vccd1 _5917_/A sky130_fd_sc_hd__xnor2_2
X_8266_ _8266_/A _8386_/B _8266_/C vssd1 vssd1 vccd1 vccd1 _8268_/B sky130_fd_sc_hd__nand3_1
X_5478_ _5478_/A _5478_/B vssd1 vssd1 vccd1 vccd1 _5484_/B sky130_fd_sc_hd__or2_1
X_7217_ _7217_/A _7217_/B vssd1 vssd1 vccd1 vccd1 _7219_/C sky130_fd_sc_hd__xnor2_1
X_4429_ _4431_/A vssd1 vssd1 vccd1 vccd1 _4429_/Y sky130_fd_sc_hd__inv_2
X_8197_ _8197_/A _8197_/B vssd1 vssd1 vccd1 vccd1 _8237_/A sky130_fd_sc_hd__xor2_1
XFILLER_59_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7148_ _6651_/A _6650_/A _6924_/A _6644_/A vssd1 vssd1 vccd1 vccd1 _7536_/B sky130_fd_sc_hd__o31a_1
XFILLER_86_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7079_ _7079_/A _7079_/B vssd1 vssd1 vccd1 vccd1 _7087_/A sky130_fd_sc_hd__xnor2_1
XFILLER_86_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4780_ _6460_/A vssd1 vssd1 vccd1 vccd1 _5335_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6450_ _8745_/Q _6450_/B vssd1 vssd1 vccd1 vccd1 _7622_/A sky130_fd_sc_hd__nand2_2
X_6381_ _6381_/A _6381_/B vssd1 vssd1 vccd1 vccd1 _6389_/B sky130_fd_sc_hd__xnor2_1
X_5401_ _8699_/Q _8700_/Q _5401_/C vssd1 vssd1 vccd1 vccd1 _5404_/B sky130_fd_sc_hd__and3_1
X_8120_ _8120_/A vssd1 vssd1 vccd1 vccd1 _8289_/B sky130_fd_sc_hd__clkbuf_2
X_5332_ _8682_/Q _5334_/B vssd1 vssd1 vccd1 vccd1 _5332_/X sky130_fd_sc_hd__or2_1
XFILLER_87_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8051_ _8051_/A _8055_/A _8051_/C vssd1 vssd1 vccd1 vccd1 _8053_/B sky130_fd_sc_hd__or3_1
X_5263_ _5263_/A _5269_/A _5263_/C _5285_/C vssd1 vssd1 vccd1 vccd1 _5263_/X sky130_fd_sc_hd__or4_1
XFILLER_68_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7002_ _7363_/B _7379_/B _7002_/C vssd1 vssd1 vccd1 vccd1 _7004_/B sky130_fd_sc_hd__or3_1
X_5194_ _5194_/A _5291_/A _4818_/A vssd1 vssd1 vccd1 vccd1 _5194_/X sky130_fd_sc_hd__or3b_1
XFILLER_68_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8953_ _8953_/A _4440_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[2] sky130_fd_sc_hd__ebufn_8
X_7904_ _7904_/A vssd1 vssd1 vccd1 vccd1 _8439_/A sky130_fd_sc_hd__clkbuf_2
X_8884_ _8884_/A _4361_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[3] sky130_fd_sc_hd__ebufn_8
XFILLER_24_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7835_ _8273_/A vssd1 vssd1 vccd1 vccd1 _8261_/A sky130_fd_sc_hd__clkbuf_2
X_7766_ _7773_/A _7766_/B vssd1 vssd1 vccd1 vccd1 _7882_/A sky130_fd_sc_hd__nand2_1
X_4978_ _4978_/A vssd1 vssd1 vccd1 vccd1 _5225_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7697_ _8325_/A _7839_/B vssd1 vssd1 vccd1 vccd1 _7712_/A sky130_fd_sc_hd__or2_1
X_6717_ _6816_/C _6717_/B vssd1 vssd1 vccd1 vccd1 _6957_/A sky130_fd_sc_hd__nand2_1
X_6648_ _6648_/A _6648_/B vssd1 vssd1 vccd1 vccd1 _6694_/A sky130_fd_sc_hd__and2_1
X_8318_ _8308_/A _8308_/B _8317_/Y vssd1 vssd1 vccd1 vccd1 _8481_/A sky130_fd_sc_hd__a21o_1
XFILLER_3_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6579_ _6570_/A _6583_/B _6571_/Y vssd1 vssd1 vccd1 vccd1 _6580_/B sky130_fd_sc_hd__a21o_1
XFILLER_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8249_ _8249_/A _8273_/B vssd1 vssd1 vccd1 vccd1 _8389_/B sky130_fd_sc_hd__nor2_2
XFILLER_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5950_ _5950_/A _5950_/B vssd1 vssd1 vccd1 vccd1 _5951_/B sky130_fd_sc_hd__or2_1
XFILLER_92_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4901_ _4901_/A _4901_/B vssd1 vssd1 vccd1 vccd1 _5100_/B sky130_fd_sc_hd__nor2_2
X_5881_ _5881_/A _5881_/B _5881_/C vssd1 vssd1 vccd1 vccd1 _5961_/B sky130_fd_sc_hd__and3_1
X_7620_ _7622_/B _7616_/X _7619_/X _7651_/B vssd1 vssd1 vccd1 vccd1 _7621_/B sky130_fd_sc_hd__a22o_1
XFILLER_21_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4832_ _4894_/B _4982_/B vssd1 vssd1 vccd1 vccd1 _5206_/A sky130_fd_sc_hd__nor2_1
X_4763_ _4897_/C vssd1 vssd1 vccd1 vccd1 _5100_/A sky130_fd_sc_hd__clkbuf_2
X_7551_ _7551_/A _7551_/B vssd1 vssd1 vccd1 vccd1 _7552_/C sky130_fd_sc_hd__xnor2_1
X_4694_ input2/X vssd1 vssd1 vccd1 vccd1 _6460_/A sky130_fd_sc_hd__buf_2
X_7482_ _7483_/B _7482_/B vssd1 vssd1 vccd1 vccd1 _7482_/X sky130_fd_sc_hd__and2b_1
X_6502_ _8737_/Q _6501_/B _6483_/X vssd1 vssd1 vccd1 vccd1 _6503_/B sky130_fd_sc_hd__o21ai_1
X_6433_ _6433_/A _6433_/B _6432_/X vssd1 vssd1 vccd1 vccd1 _6435_/B sky130_fd_sc_hd__or3b_1
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6364_ _6367_/B _6367_/C _6367_/A vssd1 vssd1 vccd1 vccd1 _6365_/C sky130_fd_sc_hd__a21oi_1
X_6295_ _6296_/A _6296_/B vssd1 vssd1 vccd1 vccd1 _6297_/A sky130_fd_sc_hd__nand2_1
X_8103_ _8103_/A _8498_/S vssd1 vssd1 vccd1 vccd1 _8121_/B sky130_fd_sc_hd__nor2_1
X_5315_ _5315_/A vssd1 vssd1 vccd1 vccd1 _5326_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_8034_ _8034_/A _8034_/B vssd1 vssd1 vccd1 vccd1 _8114_/B sky130_fd_sc_hd__xnor2_1
X_5246_ _5300_/B _5247_/B vssd1 vssd1 vccd1 vccd1 _5246_/Y sky130_fd_sc_hd__nor2_1
XFILLER_102_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5177_ _5266_/A _5283_/C _5265_/B _5066_/Y _5163_/C vssd1 vssd1 vccd1 vccd1 _5179_/C
+ sky130_fd_sc_hd__o32a_1
XFILLER_28_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8936_ _8936_/A _4424_/Y vssd1 vssd1 vccd1 vccd1 io_out[23] sky130_fd_sc_hd__ebufn_8
XFILLER_83_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7818_ _7818_/A _7924_/C vssd1 vssd1 vccd1 vccd1 _7819_/B sky130_fd_sc_hd__xnor2_1
X_7749_ _7789_/A _7789_/B vssd1 vssd1 vccd1 vccd1 _8172_/A sky130_fd_sc_hd__xnor2_4
XFILLER_61_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6080_ _6194_/A vssd1 vssd1 vccd1 vccd1 _6274_/B sky130_fd_sc_hd__clkbuf_2
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5100_ _5100_/A _5100_/B _5107_/B vssd1 vssd1 vccd1 vccd1 _5101_/B sky130_fd_sc_hd__and3_1
X_8871__88 vssd1 vssd1 vccd1 vccd1 _8871__88/HI _8980_/A sky130_fd_sc_hd__conb_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5031_ _5281_/A _5031_/B _5148_/A _5030_/Y vssd1 vssd1 vccd1 vccd1 _5031_/X sky130_fd_sc_hd__or4b_1
XFILLER_97_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6982_ _6982_/A _6982_/B vssd1 vssd1 vccd1 vccd1 _6984_/A sky130_fd_sc_hd__xnor2_1
XFILLER_25_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8721_ _8765_/CLK _8721_/D vssd1 vssd1 vccd1 vccd1 _8721_/Q sky130_fd_sc_hd__dfxtp_1
X_5933_ _5933_/A _6302_/A vssd1 vssd1 vccd1 vccd1 _5934_/B sky130_fd_sc_hd__xnor2_1
X_5864_ _5864_/A _5864_/B vssd1 vssd1 vccd1 vccd1 _5864_/Y sky130_fd_sc_hd__nand2_1
X_8652_ _8778_/CLK _8652_/D vssd1 vssd1 vccd1 vccd1 _8652_/Q sky130_fd_sc_hd__dfxtp_1
X_8583_ _8586_/B _8582_/Y _8578_/A _8578_/B vssd1 vssd1 vccd1 vccd1 _8583_/X sky130_fd_sc_hd__a211o_1
X_7603_ _8783_/Q vssd1 vssd1 vccd1 vccd1 _8626_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4815_ _4767_/B _4813_/X _4814_/Y _5315_/A _4814_/A vssd1 vssd1 vccd1 vccd1 _4816_/B
+ sky130_fd_sc_hd__a32o_1
X_5795_ _5792_/X _5793_/Y _5714_/X _5715_/Y vssd1 vssd1 vccd1 vccd1 _5801_/B sky130_fd_sc_hd__o211a_1
X_7534_ _7534_/A _7540_/A _7540_/B _7540_/C vssd1 vssd1 vccd1 vccd1 _7552_/B sky130_fd_sc_hd__or4_1
X_4746_ _4771_/A _5259_/D _4741_/A _5249_/B vssd1 vssd1 vccd1 vccd1 _4747_/C sky130_fd_sc_hd__a31o_1
X_4677_ _8650_/Q _4678_/B vssd1 vssd1 vccd1 vccd1 _4679_/B sky130_fd_sc_hd__or2_1
X_7465_ _7465_/A _7465_/B _7465_/C vssd1 vssd1 vccd1 vccd1 _7467_/A sky130_fd_sc_hd__and3_1
X_6416_ _6416_/A _6416_/B vssd1 vssd1 vccd1 vccd1 _6423_/B sky130_fd_sc_hd__and2_1
X_7396_ _7396_/A _7446_/A vssd1 vssd1 vccd1 vccd1 _7399_/A sky130_fd_sc_hd__xor2_2
X_6347_ _6284_/A _6345_/X _6346_/X vssd1 vssd1 vccd1 vccd1 _6348_/B sky130_fd_sc_hd__o21a_1
XFILLER_103_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6278_ _6278_/A _6278_/B vssd1 vssd1 vccd1 vccd1 _6279_/B sky130_fd_sc_hd__nor2_1
XFILLER_102_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8017_ _8060_/B _8016_/C _8016_/A vssd1 vssd1 vccd1 vccd1 _8018_/C sky130_fd_sc_hd__a21o_1
X_5229_ _5047_/A _5234_/A _5069_/D _5228_/X vssd1 vssd1 vccd1 vccd1 _5229_/Y sky130_fd_sc_hd__a211oi_1
XFILLER_48_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8919_ _8919_/A _4404_/Y vssd1 vssd1 vccd1 vccd1 io_out[6] sky130_fd_sc_hd__ebufn_8
XFILLER_72_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_2_3_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_79_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4600_ _4600_/A vssd1 vssd1 vccd1 vccd1 _8933_/A sky130_fd_sc_hd__clkbuf_2
X_5580_ _5979_/A _5687_/A vssd1 vssd1 vccd1 vccd1 _5749_/A sky130_fd_sc_hd__nand2_2
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4531_ _8663_/Q vssd1 vssd1 vccd1 vccd1 _4774_/A sky130_fd_sc_hd__clkbuf_1
X_4462_ _4462_/A vssd1 vssd1 vccd1 vccd1 _4462_/Y sky130_fd_sc_hd__inv_2
X_7250_ _7525_/A _7528_/B _7525_/C _7533_/A _7249_/X vssd1 vssd1 vccd1 vccd1 _7524_/S
+ sky130_fd_sc_hd__a41o_1
X_6201_ _6277_/B _6277_/C vssd1 vssd1 vccd1 vccd1 _6278_/B sky130_fd_sc_hd__xnor2_1
XFILLER_98_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4393_ _4394_/A vssd1 vssd1 vccd1 vccd1 _4393_/Y sky130_fd_sc_hd__inv_2
X_7181_ _7182_/A _7181_/B vssd1 vssd1 vccd1 vccd1 _7285_/B sky130_fd_sc_hd__nor2_1
X_6132_ _6132_/A _6132_/B vssd1 vssd1 vccd1 vccd1 _6365_/B sky130_fd_sc_hd__nor2_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6063_ _6178_/A _6063_/B vssd1 vssd1 vccd1 vccd1 _6064_/B sky130_fd_sc_hd__nor2_1
XFILLER_85_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5014_ _5006_/X _5012_/X _5286_/A _4891_/B vssd1 vssd1 vccd1 vccd1 _5014_/X sky130_fd_sc_hd__a211o_1
XFILLER_38_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6965_ _6965_/A _6965_/B vssd1 vssd1 vccd1 vccd1 _7080_/D sky130_fd_sc_hd__xnor2_2
X_5916_ _5916_/A _5916_/B vssd1 vssd1 vccd1 vccd1 _6059_/A sky130_fd_sc_hd__nand2_1
XFILLER_81_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8704_ _8704_/CLK _8704_/D vssd1 vssd1 vccd1 vccd1 _8704_/Q sky130_fd_sc_hd__dfxtp_1
X_6896_ _6879_/A _6879_/B _6861_/A vssd1 vssd1 vccd1 vccd1 _6920_/A sky130_fd_sc_hd__a21o_1
X_8635_ _8730_/CLK _8635_/D vssd1 vssd1 vccd1 vccd1 _8635_/Q sky130_fd_sc_hd__dfxtp_1
X_5847_ _5847_/A _5887_/B _5847_/C vssd1 vssd1 vccd1 vccd1 _5886_/A sky130_fd_sc_hd__and3_1
X_5778_ _5783_/A _5851_/C vssd1 vssd1 vccd1 vccd1 _5849_/B sky130_fd_sc_hd__xnor2_1
X_8566_ _8567_/A _8567_/B vssd1 vssd1 vccd1 vccd1 _8571_/A sky130_fd_sc_hd__nand2_1
X_8497_ _8497_/A _8497_/B vssd1 vssd1 vccd1 vccd1 _8499_/A sky130_fd_sc_hd__or2_1
X_7517_ _7538_/A _7537_/A vssd1 vssd1 vccd1 vccd1 _7518_/B sky130_fd_sc_hd__or2_1
X_4729_ _4818_/A _4818_/B vssd1 vssd1 vccd1 vccd1 _5170_/A sky130_fd_sc_hd__or2_2
X_7448_ _7489_/A _7489_/B vssd1 vssd1 vccd1 vccd1 _7449_/B sky130_fd_sc_hd__nand2_1
XFILLER_101_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7379_ _7391_/B _7379_/B vssd1 vssd1 vccd1 vccd1 _7489_/B sky130_fd_sc_hd__nor2_2
XFILLER_76_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8841__58 vssd1 vssd1 vccd1 vccd1 _8841__58/HI _8950_/A sky130_fd_sc_hd__conb_1
XFILLER_63_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6750_ _8754_/Q _7842_/B vssd1 vssd1 vccd1 vccd1 _6752_/A sky130_fd_sc_hd__nor2_1
X_5701_ _5991_/A _5701_/B vssd1 vssd1 vccd1 vccd1 _5702_/B sky130_fd_sc_hd__and2_1
XFILLER_16_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6681_ _7229_/A vssd1 vssd1 vccd1 vccd1 _7181_/B sky130_fd_sc_hd__buf_2
XFILLER_31_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8420_ _8420_/A _8420_/B vssd1 vssd1 vccd1 vccd1 _8494_/B sky130_fd_sc_hd__xnor2_1
X_5632_ _5632_/A vssd1 vssd1 vccd1 vccd1 _5824_/B sky130_fd_sc_hd__clkbuf_2
X_8351_ _8418_/A _8351_/B vssd1 vssd1 vccd1 vccd1 _8360_/A sky130_fd_sc_hd__xnor2_1
X_5563_ _6615_/B _6409_/A vssd1 vssd1 vccd1 vccd1 _5564_/B sky130_fd_sc_hd__and2b_1
X_4514_ _8669_/Q vssd1 vssd1 vccd1 vccd1 _7700_/A sky130_fd_sc_hd__buf_2
X_7302_ _7302_/A _7302_/B vssd1 vssd1 vccd1 vccd1 _7377_/A sky130_fd_sc_hd__nor2_2
X_8282_ _8282_/A _8281_/X vssd1 vssd1 vccd1 vccd1 _8364_/B sky130_fd_sc_hd__or2b_1
X_5494_ _5494_/A _6621_/B vssd1 vssd1 vccd1 vccd1 _5552_/B sky130_fd_sc_hd__nand2_1
XFILLER_104_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4445_ _4457_/A vssd1 vssd1 vccd1 vccd1 _4450_/A sky130_fd_sc_hd__buf_4
X_7233_ _7327_/B _7233_/B vssd1 vssd1 vccd1 vccd1 _7336_/B sky130_fd_sc_hd__xnor2_1
X_4376_ _4376_/A vssd1 vssd1 vccd1 vccd1 _4376_/Y sky130_fd_sc_hd__inv_2
X_7164_ _7060_/A _7060_/B _7163_/X vssd1 vssd1 vccd1 vccd1 _7242_/A sky130_fd_sc_hd__a21o_1
X_6115_ _6116_/A _6116_/B vssd1 vssd1 vccd1 vccd1 _6162_/A sky130_fd_sc_hd__nor2_1
XFILLER_98_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7095_ _7097_/B _7097_/A vssd1 vssd1 vccd1 vccd1 _7096_/C sky130_fd_sc_hd__or2b_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6046_ _6050_/A _6050_/B vssd1 vssd1 vccd1 vccd1 _6047_/B sky130_fd_sc_hd__xor2_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7997_ _8172_/B vssd1 vssd1 vccd1 vccd1 _8273_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_54_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6948_ _6949_/A _6949_/B vssd1 vssd1 vccd1 vccd1 _6948_/Y sky130_fd_sc_hd__nand2_1
X_6879_ _6879_/A _6879_/B vssd1 vssd1 vccd1 vccd1 _6894_/B sky130_fd_sc_hd__xnor2_1
X_8618_ _8626_/A _8609_/A _8617_/X _7642_/X vssd1 vssd1 vccd1 vccd1 _8783_/D sky130_fd_sc_hd__o211a_1
XFILLER_10_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8549_ _8549_/A _8549_/B _8549_/C vssd1 vssd1 vccd1 vccd1 _8549_/X sky130_fd_sc_hd__and3_1
XFILLER_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7920_ _7919_/A _7919_/B _7919_/C vssd1 vssd1 vccd1 vccd1 _7921_/C sky130_fd_sc_hd__a21o_1
XFILLER_36_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7851_ _7938_/A _7938_/B vssd1 vssd1 vccd1 vccd1 _7959_/A sky130_fd_sc_hd__xnor2_1
X_6802_ _6802_/A _6802_/B vssd1 vssd1 vccd1 vccd1 _6804_/B sky130_fd_sc_hd__nand2_1
XFILLER_90_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7782_ _8025_/A _8354_/A vssd1 vssd1 vccd1 vccd1 _7783_/B sky130_fd_sc_hd__nor2_1
X_4994_ _5155_/C _5050_/D _4991_/Y _4993_/Y vssd1 vssd1 vccd1 vccd1 _4995_/D sky130_fd_sc_hd__o31a_1
X_6733_ _7685_/A _8751_/Q vssd1 vssd1 vccd1 vccd1 _6735_/A sky130_fd_sc_hd__and2b_1
X_6664_ _7587_/A _6673_/B vssd1 vssd1 vccd1 vccd1 _7363_/A sky130_fd_sc_hd__and2_1
X_8403_ _8403_/A _8403_/B vssd1 vssd1 vccd1 vccd1 _8404_/B sky130_fd_sc_hd__xnor2_1
X_5615_ _5615_/A _5615_/B vssd1 vssd1 vccd1 vccd1 _5615_/X sky130_fd_sc_hd__or2_1
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6595_ _6758_/A _8747_/Q vssd1 vssd1 vccd1 vccd1 _6602_/B sky130_fd_sc_hd__nand2_1
X_8334_ _8414_/A _8414_/B vssd1 vssd1 vccd1 vccd1 _8335_/B sky130_fd_sc_hd__xor2_1
X_5546_ _5655_/B vssd1 vssd1 vccd1 vccd1 _6166_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_3_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8265_ _8264_/B _8386_/A _8264_/A vssd1 vssd1 vccd1 vccd1 _8266_/C sky130_fd_sc_hd__a21o_1
X_5477_ _5478_/A _5477_/B vssd1 vssd1 vccd1 vccd1 _5480_/C sky130_fd_sc_hd__nand2_1
X_4428_ _4431_/A vssd1 vssd1 vccd1 vccd1 _4428_/Y sky130_fd_sc_hd__inv_2
X_7216_ _7216_/A _7216_/B vssd1 vssd1 vccd1 vccd1 _7217_/B sky130_fd_sc_hd__xor2_1
X_8196_ _8122_/Y _8358_/A _8336_/A _8195_/Y vssd1 vssd1 vccd1 vccd1 _8197_/B sky130_fd_sc_hd__o31a_1
XFILLER_98_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7147_ _7147_/A _7147_/B vssd1 vssd1 vccd1 vccd1 _7536_/A sky130_fd_sc_hd__xnor2_1
X_4359_ _4363_/A vssd1 vssd1 vccd1 vccd1 _4359_/Y sky130_fd_sc_hd__inv_2
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7078_ _7078_/A _7078_/B vssd1 vssd1 vccd1 vccd1 _7082_/A sky130_fd_sc_hd__nand2_1
XFILLER_48_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6029_ _6029_/A _6029_/B vssd1 vssd1 vccd1 vccd1 _6030_/B sky130_fd_sc_hd__xor2_1
XFILLER_46_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8811__28 vssd1 vssd1 vccd1 vccd1 _8811__28/HI _8906_/A sky130_fd_sc_hd__conb_1
XFILLER_64_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6380_ _6390_/A _6390_/B _6388_/B vssd1 vssd1 vccd1 vccd1 _6380_/X sky130_fd_sc_hd__or3_1
X_5400_ _5400_/A _5400_/B vssd1 vssd1 vccd1 vccd1 _8699_/D sky130_fd_sc_hd__nor2_1
X_5331_ _8756_/Q _5320_/X _5330_/X _5324_/X vssd1 vssd1 vccd1 vccd1 _8681_/D sky130_fd_sc_hd__o211a_1
X_8050_ _8057_/B _8048_/X _7972_/A _7974_/A vssd1 vssd1 vccd1 vccd1 _8051_/C sky130_fd_sc_hd__a211oi_1
X_7001_ _7001_/A _6904_/B vssd1 vssd1 vccd1 vccd1 _7169_/A sky130_fd_sc_hd__or2b_1
X_5262_ _5009_/C _5107_/A _5135_/B vssd1 vssd1 vccd1 vccd1 _5285_/C sky130_fd_sc_hd__a21o_1
XFILLER_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5193_ _5179_/B _5291_/C _5186_/X _5192_/X vssd1 vssd1 vccd1 vccd1 _5194_/A sky130_fd_sc_hd__o31a_1
XFILLER_68_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8952_ _8952_/A _4442_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[1] sky130_fd_sc_hd__ebufn_8
XFILLER_83_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7903_ _7903_/A vssd1 vssd1 vccd1 vccd1 _8008_/A sky130_fd_sc_hd__clkbuf_2
X_8883_ _8883_/A _4360_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[2] sky130_fd_sc_hd__ebufn_8
X_7834_ _7834_/A _7894_/B vssd1 vssd1 vccd1 vccd1 _7892_/A sky130_fd_sc_hd__xor2_1
X_7765_ _7940_/A _7712_/A _8332_/C _7764_/Y _7715_/X vssd1 vssd1 vccd1 vccd1 _7766_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_51_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4977_ _4977_/A vssd1 vssd1 vccd1 vccd1 _4977_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6716_ _6810_/A _7302_/B _7205_/B _7030_/A vssd1 vssd1 vccd1 vccd1 _6717_/B sky130_fd_sc_hd__o22ai_1
X_7696_ _7696_/A vssd1 vssd1 vccd1 vccd1 _7839_/B sky130_fd_sc_hd__clkbuf_2
X_6647_ _7123_/A _6647_/B vssd1 vssd1 vccd1 vccd1 _6650_/A sky130_fd_sc_hd__nor2_1
X_6578_ _6578_/A _6578_/B vssd1 vssd1 vccd1 vccd1 _6580_/A sky130_fd_sc_hd__nor2_1
X_8877__94 vssd1 vssd1 vccd1 vccd1 _8877__94/HI _8986_/A sky130_fd_sc_hd__conb_1
X_5529_ _5922_/A _6107_/A _5528_/Y vssd1 vssd1 vccd1 vccd1 _5532_/A sky130_fd_sc_hd__a21oi_1
X_8317_ _8317_/A _8317_/B vssd1 vssd1 vccd1 vccd1 _8317_/Y sky130_fd_sc_hd__nor2_1
XFILLER_59_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8248_ _8450_/A _8248_/B _8248_/C vssd1 vssd1 vccd1 vccd1 _8254_/A sky130_fd_sc_hd__and3_1
X_8179_ _8179_/A _8179_/B vssd1 vssd1 vccd1 vccd1 _8246_/B sky130_fd_sc_hd__xnor2_2
XFILLER_78_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5880_ _5883_/A _5879_/C _5879_/A vssd1 vssd1 vccd1 vccd1 _5881_/C sky130_fd_sc_hd__o21ai_1
XFILLER_73_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4900_ _5083_/B _4912_/B vssd1 vssd1 vccd1 vccd1 _5288_/C sky130_fd_sc_hd__nor2_1
X_4831_ _4925_/B vssd1 vssd1 vccd1 vccd1 _4982_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_60_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4762_ _4762_/A vssd1 vssd1 vccd1 vccd1 _4897_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7550_ _7541_/X _7549_/X _5491_/X _8757_/Q vssd1 vssd1 vccd1 vccd1 _8757_/D sky130_fd_sc_hd__o2bb2a_1
X_4693_ _5136_/A _4771_/A vssd1 vssd1 vccd1 vccd1 _4732_/B sky130_fd_sc_hd__nand2_1
X_7481_ _7481_/A _7481_/B vssd1 vssd1 vccd1 vccd1 _7503_/A sky130_fd_sc_hd__xnor2_1
X_6501_ _8737_/Q _6501_/B vssd1 vssd1 vccd1 vccd1 _6506_/C sky130_fd_sc_hd__and2_1
X_6432_ _6428_/A _6431_/X _6432_/S vssd1 vssd1 vccd1 vccd1 _6432_/X sky130_fd_sc_hd__mux2_1
X_6363_ _6363_/A _6363_/B vssd1 vssd1 vccd1 vccd1 _6365_/A sky130_fd_sc_hd__xor2_1
X_8102_ _8102_/A _8102_/B vssd1 vssd1 vccd1 vccd1 _8498_/S sky130_fd_sc_hd__nand2_1
X_6294_ _6294_/A _6294_/B vssd1 vssd1 vccd1 vccd1 _6296_/B sky130_fd_sc_hd__xor2_1
XFILLER_88_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5314_ _8716_/Q _5307_/X _5313_/X _5311_/X vssd1 vssd1 vccd1 vccd1 _8674_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8033_ _8099_/A _8293_/A vssd1 vssd1 vccd1 vccd1 _8034_/B sky130_fd_sc_hd__nor2_1
X_5245_ _4977_/A _5196_/X _5244_/X _5296_/A vssd1 vssd1 vccd1 vccd1 _5245_/Y sky130_fd_sc_hd__o211ai_1
X_5176_ _5176_/A _5281_/A _5283_/C _5178_/B vssd1 vssd1 vccd1 vccd1 _5176_/X sky130_fd_sc_hd__or4_1
XFILLER_56_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8935_ _8935_/A _4423_/Y vssd1 vssd1 vccd1 vccd1 io_out[22] sky130_fd_sc_hd__ebufn_8
XFILLER_83_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_3_5_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
X_7817_ _7998_/A _8010_/A _7816_/X vssd1 vssd1 vccd1 vccd1 _7924_/C sky130_fd_sc_hd__o21a_1
X_7748_ _7788_/A _7788_/B _7725_/A vssd1 vssd1 vccd1 vccd1 _7789_/A sky130_fd_sc_hd__a21o_2
X_7679_ _7679_/A _8770_/Q vssd1 vssd1 vccd1 vccd1 _7688_/A sky130_fd_sc_hd__or2b_2
XFILLER_3_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5030_ _5250_/D _5211_/A _5128_/A vssd1 vssd1 vccd1 vccd1 _5030_/Y sky130_fd_sc_hd__nor3_1
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6981_ _7075_/A _7075_/B _6978_/B _7070_/A _7070_/B vssd1 vssd1 vccd1 vccd1 _6983_/A
+ sky130_fd_sc_hd__a32o_1
X_5932_ _5932_/A _6016_/A vssd1 vssd1 vccd1 vccd1 _6302_/A sky130_fd_sc_hd__xnor2_4
XFILLER_65_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8720_ _8720_/CLK _8720_/D vssd1 vssd1 vccd1 vccd1 _8720_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5863_ _5937_/A _5937_/B vssd1 vssd1 vccd1 vccd1 _5942_/A sky130_fd_sc_hd__xnor2_1
X_8651_ _8723_/CLK _8651_/D vssd1 vssd1 vccd1 vccd1 _8651_/Q sky130_fd_sc_hd__dfxtp_1
X_5794_ _5714_/X _5715_/Y _5792_/X _5793_/Y vssd1 vssd1 vccd1 vccd1 _5801_/A sky130_fd_sc_hd__a211oi_2
X_8582_ _8582_/A _8582_/B vssd1 vssd1 vccd1 vccd1 _8582_/Y sky130_fd_sc_hd__nand2_1
X_7602_ _7602_/A _7619_/B _7619_/C _7602_/D vssd1 vssd1 vccd1 vccd1 _7602_/X sky130_fd_sc_hd__or4_1
XFILLER_33_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4814_ _4814_/A _4814_/B _4814_/C _4814_/D vssd1 vssd1 vccd1 vccd1 _4814_/Y sky130_fd_sc_hd__nand4_1
X_4745_ _4745_/A _5247_/B vssd1 vssd1 vccd1 vccd1 _4751_/B sky130_fd_sc_hd__nor2_1
X_7533_ _7533_/A _7533_/B vssd1 vssd1 vccd1 vccd1 _7540_/C sky130_fd_sc_hd__xor2_2
XFILLER_21_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7464_ _7395_/A _7395_/B _7463_/X vssd1 vssd1 vccd1 vccd1 _7465_/C sky130_fd_sc_hd__a21oi_1
X_4676_ _4678_/B _4676_/B vssd1 vssd1 vccd1 vccd1 _8649_/D sky130_fd_sc_hd__nor2_1
X_6415_ _6415_/A _6415_/B vssd1 vssd1 vccd1 vccd1 _6416_/B sky130_fd_sc_hd__or2_1
X_7395_ _7395_/A _7395_/B vssd1 vssd1 vccd1 vccd1 _7446_/A sky130_fd_sc_hd__xnor2_2
X_6346_ _6346_/A _6283_/B vssd1 vssd1 vccd1 vccd1 _6346_/X sky130_fd_sc_hd__or2b_1
X_8847__64 vssd1 vssd1 vccd1 vccd1 _8847__64/HI _8956_/A sky130_fd_sc_hd__conb_1
XFILLER_103_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8016_ _8016_/A _8060_/B _8016_/C vssd1 vssd1 vccd1 vccd1 _8059_/A sky130_fd_sc_hd__nand3_1
X_6277_ _6278_/A _6277_/B _6277_/C vssd1 vssd1 vccd1 vccd1 _6279_/A sky130_fd_sc_hd__and3_1
XFILLER_69_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5228_ _5228_/A _5228_/B _5228_/C vssd1 vssd1 vccd1 vccd1 _5228_/X sky130_fd_sc_hd__or3_1
X_5159_ _5263_/A _5159_/B _5278_/B _5159_/D vssd1 vssd1 vccd1 vccd1 _5159_/X sky130_fd_sc_hd__or4_1
XFILLER_56_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8918_ _8918_/A _4403_/Y vssd1 vssd1 vccd1 vccd1 io_out[5] sky130_fd_sc_hd__ebufn_8
XFILLER_72_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4530_ _4804_/A _5298_/A _4870_/A vssd1 vssd1 vccd1 vccd1 _4568_/B sky130_fd_sc_hd__nand3_1
X_4461_ _4462_/A vssd1 vssd1 vccd1 vccd1 _4461_/Y sky130_fd_sc_hd__inv_2
X_6200_ _6200_/A _6200_/B vssd1 vssd1 vccd1 vccd1 _6277_/C sky130_fd_sc_hd__xnor2_1
X_7180_ _7318_/B _7180_/B vssd1 vssd1 vccd1 vccd1 _7194_/A sky130_fd_sc_hd__nand2_1
X_6131_ _6367_/B _6367_/C _6127_/Y _6367_/A vssd1 vssd1 vccd1 vccd1 _6360_/B sky130_fd_sc_hd__a211o_1
X_4392_ _4394_/A vssd1 vssd1 vccd1 vccd1 _4392_/Y sky130_fd_sc_hd__inv_2
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6062_ _6252_/A _6062_/B vssd1 vssd1 vccd1 vccd1 _6063_/B sky130_fd_sc_hd__and2_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5013_ _5138_/A _5251_/A vssd1 vssd1 vccd1 vccd1 _5286_/A sky130_fd_sc_hd__or2_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6964_ _7118_/A _7123_/B vssd1 vssd1 vccd1 vccd1 _6965_/B sky130_fd_sc_hd__nand2_1
X_5915_ _6169_/B vssd1 vssd1 vccd1 vccd1 _6171_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_81_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6895_ _6889_/A _6889_/B _6894_/X vssd1 vssd1 vccd1 vccd1 _6941_/A sky130_fd_sc_hd__o21a_1
X_8703_ _8704_/CLK _8703_/D vssd1 vssd1 vccd1 vccd1 _8703_/Q sky130_fd_sc_hd__dfxtp_1
X_5846_ _5887_/A _5845_/C _5845_/A vssd1 vssd1 vccd1 vccd1 _5847_/C sky130_fd_sc_hd__a21o_1
XFILLER_34_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8634_ _8732_/CLK _8634_/D vssd1 vssd1 vccd1 vccd1 _8634_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5777_ _5872_/A _5777_/B vssd1 vssd1 vccd1 vccd1 _5851_/C sky130_fd_sc_hd__nor2_2
X_8565_ _8565_/A _8565_/B _8565_/C _8565_/D vssd1 vssd1 vccd1 vccd1 _8578_/B sky130_fd_sc_hd__or4_4
X_8496_ _8358_/B _8356_/B _8496_/S vssd1 vssd1 vccd1 vccd1 _8497_/B sky130_fd_sc_hd__mux2_1
XFILLER_21_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7516_ _7516_/A _7516_/B vssd1 vssd1 vccd1 vccd1 _7551_/A sky130_fd_sc_hd__or2_1
X_4728_ _4734_/B vssd1 vssd1 vccd1 vccd1 _4818_/B sky130_fd_sc_hd__clkbuf_2
X_4659_ _8644_/Q _4661_/C _4679_/A vssd1 vssd1 vccd1 vccd1 _4659_/Y sky130_fd_sc_hd__o21ai_1
X_7447_ _7399_/A _7399_/B _7446_/X vssd1 vssd1 vccd1 vccd1 _7455_/A sky130_fd_sc_hd__o21ai_1
XFILLER_103_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7378_ _7378_/A _7388_/S vssd1 vssd1 vccd1 vccd1 _7384_/A sky130_fd_sc_hd__nand2_1
X_6329_ _6192_/A _6274_/Y _5827_/X vssd1 vssd1 vccd1 vccd1 _6330_/B sky130_fd_sc_hd__o21ba_1
XFILLER_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5700_ _5700_/A _5926_/A _5700_/C vssd1 vssd1 vccd1 vccd1 _6377_/A sky130_fd_sc_hd__and3_1
XFILLER_16_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6680_ _7363_/B _7379_/B _6688_/A vssd1 vssd1 vccd1 vccd1 _7229_/A sky130_fd_sc_hd__or3_2
X_5631_ _6092_/A vssd1 vssd1 vccd1 vccd1 _6197_/A sky130_fd_sc_hd__buf_2
X_8350_ _8098_/A _8357_/A _8349_/X vssd1 vssd1 vccd1 vccd1 _8351_/B sky130_fd_sc_hd__o21a_1
X_5562_ _8720_/Q _8657_/Q vssd1 vssd1 vccd1 vccd1 _5564_/A sky130_fd_sc_hd__and2b_1
X_8281_ _8280_/A _8280_/B _8280_/C _8280_/D vssd1 vssd1 vccd1 vccd1 _8281_/X sky130_fd_sc_hd__a22o_1
X_7301_ _7301_/A _7309_/B vssd1 vssd1 vccd1 vccd1 _7305_/A sky130_fd_sc_hd__nand2_1
X_4513_ _4778_/A vssd1 vssd1 vccd1 vccd1 _4549_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5493_ _5493_/A vssd1 vssd1 vccd1 vccd1 _5552_/A sky130_fd_sc_hd__clkbuf_4
X_7232_ _7392_/B _7181_/B _7230_/A _7052_/B vssd1 vssd1 vccd1 vccd1 _7233_/B sky130_fd_sc_hd__o22a_1
X_4444_ _4444_/A vssd1 vssd1 vccd1 vccd1 _4444_/Y sky130_fd_sc_hd__clkinv_2
X_8817__34 vssd1 vssd1 vccd1 vccd1 _8817__34/HI _8912_/A sky130_fd_sc_hd__conb_1
X_4375_ _4376_/A vssd1 vssd1 vccd1 vccd1 _4375_/Y sky130_fd_sc_hd__inv_2
X_7163_ _7059_/B _7163_/B vssd1 vssd1 vccd1 vccd1 _7163_/X sky130_fd_sc_hd__and2b_1
X_6114_ _5946_/B _6038_/B _6036_/Y vssd1 vssd1 vccd1 vccd1 _6116_/B sky130_fd_sc_hd__a21o_1
X_7094_ _6834_/B _6691_/B _6693_/B _6814_/A vssd1 vssd1 vccd1 vccd1 _7097_/A sky130_fd_sc_hd__a22o_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6045_ _6045_/A _6045_/B vssd1 vssd1 vccd1 vccd1 _6050_/B sky130_fd_sc_hd__xnor2_1
XFILLER_100_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7996_ _7996_/A _8158_/A vssd1 vssd1 vccd1 vccd1 _8001_/A sky130_fd_sc_hd__nand2_1
X_6947_ _7181_/B _6947_/B vssd1 vssd1 vccd1 vccd1 _6949_/B sky130_fd_sc_hd__nand2_1
X_6878_ _6922_/A _6922_/B vssd1 vssd1 vccd1 vccd1 _6879_/B sky130_fd_sc_hd__xor2_1
XFILLER_22_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5829_ _5829_/A _5829_/B vssd1 vssd1 vccd1 vccd1 _5830_/C sky130_fd_sc_hd__xnor2_1
X_8617_ _8627_/S _8616_/Y _8603_/A vssd1 vssd1 vccd1 vccd1 _8617_/X sky130_fd_sc_hd__a21o_1
X_8548_ _8549_/B _8549_/C _8549_/A vssd1 vssd1 vccd1 vccd1 _8548_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_22_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8479_ _8479_/A _8479_/B vssd1 vssd1 vccd1 vccd1 _8550_/B sky130_fd_sc_hd__xor2_1
XFILLER_78_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7850_ _7854_/B _7850_/B vssd1 vssd1 vccd1 vccd1 _7938_/B sky130_fd_sc_hd__xnor2_1
XFILLER_63_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6801_ _6801_/A _6801_/B _6801_/C vssd1 vssd1 vccd1 vccd1 _6802_/B sky130_fd_sc_hd__nand3_1
XFILLER_90_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7781_ _8568_/A _8348_/A vssd1 vssd1 vccd1 vccd1 _7784_/A sky130_fd_sc_hd__nor2_1
X_4993_ _4947_/A _4982_/B _4985_/Y _4964_/X _5176_/A vssd1 vssd1 vccd1 vccd1 _4993_/Y
+ sky130_fd_sc_hd__o221ai_1
X_6732_ _8669_/Q _8752_/Q vssd1 vssd1 vccd1 vccd1 _6732_/X sky130_fd_sc_hd__or2b_1
X_6663_ _6696_/A _6702_/A _6695_/B _6657_/A _6662_/X vssd1 vssd1 vccd1 vccd1 _6674_/D
+ sky130_fd_sc_hd__a311o_2
X_8402_ _8402_/A _8411_/B vssd1 vssd1 vccd1 vccd1 _8403_/B sky130_fd_sc_hd__xnor2_1
X_5614_ _6068_/A _5727_/A vssd1 vssd1 vccd1 vccd1 _5625_/A sky130_fd_sc_hd__nand2_1
X_6594_ _6569_/A _6602_/A _6591_/X _6593_/X vssd1 vssd1 vccd1 vccd1 _8752_/D sky130_fd_sc_hd__a31o_1
X_8333_ _8497_/A _8333_/B _8417_/B vssd1 vssd1 vccd1 vccd1 _8414_/B sky130_fd_sc_hd__and3b_1
X_5545_ _5554_/A _5554_/B vssd1 vssd1 vccd1 vccd1 _5655_/B sky130_fd_sc_hd__xor2_2
X_8264_ _8264_/A _8264_/B _8386_/A vssd1 vssd1 vccd1 vccd1 _8386_/B sky130_fd_sc_hd__nand3_1
X_5476_ _5450_/A _5474_/X _5485_/S _5449_/X _5484_/A vssd1 vssd1 vccd1 vccd1 _8711_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_2_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4427_ _4431_/A vssd1 vssd1 vccd1 vccd1 _4427_/Y sky130_fd_sc_hd__inv_2
X_8195_ _8122_/Y _8348_/A _8194_/B vssd1 vssd1 vccd1 vccd1 _8195_/Y sky130_fd_sc_hd__o21ai_1
X_7215_ _7325_/B _7215_/B vssd1 vssd1 vccd1 vccd1 _7216_/B sky130_fd_sc_hd__xnor2_1
X_7146_ _7146_/A _7146_/B vssd1 vssd1 vccd1 vccd1 _7538_/A sky130_fd_sc_hd__xnor2_1
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4358_ _4489_/A vssd1 vssd1 vccd1 vccd1 _4363_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7077_ _7105_/A _7105_/B vssd1 vssd1 vccd1 vccd1 _7078_/A sky130_fd_sc_hd__nand2_1
X_6028_ _6119_/B _6028_/B vssd1 vssd1 vccd1 vccd1 _6029_/B sky130_fd_sc_hd__nor2_1
XFILLER_27_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7979_ _8139_/B _7979_/B vssd1 vssd1 vccd1 vccd1 _7979_/X sky130_fd_sc_hd__xor2_1
XFILLER_54_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5330_ _8681_/Q _5334_/B vssd1 vssd1 vccd1 vccd1 _5330_/X sky130_fd_sc_hd__or2_1
Xclkbuf_4_7_0_wb_clk_i clkbuf_4_7_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _8720_/CLK
+ sky130_fd_sc_hd__clkbuf_2
X_5261_ _5283_/B _5261_/B _5291_/A _5261_/D vssd1 vssd1 vccd1 vccd1 _5261_/X sky130_fd_sc_hd__or4_1
X_7000_ _7000_/A _7000_/B vssd1 vssd1 vccd1 vccd1 _7025_/A sky130_fd_sc_hd__nand2_1
X_5192_ _5192_/A _5192_/B _5265_/C _5192_/D vssd1 vssd1 vccd1 vccd1 _5192_/X sky130_fd_sc_hd__or4_1
XFILLER_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8951_ _8951_/A _4486_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[0] sky130_fd_sc_hd__ebufn_8
X_7902_ _7902_/A _7902_/B _8155_/C vssd1 vssd1 vccd1 vccd1 _7903_/A sky130_fd_sc_hd__and3_1
XFILLER_24_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8882_ _8882_/A _4359_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[1] sky130_fd_sc_hd__ebufn_8
X_7833_ _8568_/D _8165_/B _7833_/C vssd1 vssd1 vccd1 vccd1 _7894_/B sky130_fd_sc_hd__and3_1
X_7764_ _7764_/A _7764_/B vssd1 vssd1 vccd1 vccd1 _7764_/Y sky130_fd_sc_hd__nand2_1
XFILLER_51_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6715_ _7302_/B _7205_/B _6725_/B vssd1 vssd1 vccd1 vccd1 _6816_/C sky130_fd_sc_hd__or3_1
X_4976_ _5249_/B _4741_/A _5247_/B vssd1 vssd1 vccd1 vccd1 _4977_/A sky130_fd_sc_hd__o21a_1
X_7695_ _7762_/A _7708_/B vssd1 vssd1 vccd1 vccd1 _7696_/A sky130_fd_sc_hd__xor2_1
X_6646_ _6646_/A vssd1 vssd1 vccd1 vccd1 _7123_/A sky130_fd_sc_hd__clkbuf_2
X_6577_ _6577_/A _8747_/Q vssd1 vssd1 vccd1 vccd1 _6578_/B sky130_fd_sc_hd__nor2_1
X_5528_ _6378_/A _5531_/D vssd1 vssd1 vccd1 vccd1 _5528_/Y sky130_fd_sc_hd__nor2_1
X_8316_ _8552_/A _8554_/B _8552_/B vssd1 vssd1 vccd1 vccd1 _8549_/C sky130_fd_sc_hd__o21ai_1
X_8247_ _8187_/A _8187_/B _8246_/X vssd1 vssd1 vccd1 vccd1 _8285_/A sky130_fd_sc_hd__a21oi_2
X_5459_ _5494_/A _5454_/B _5453_/A vssd1 vssd1 vccd1 vccd1 _5460_/B sky130_fd_sc_hd__o21a_1
XFILLER_59_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8178_ _8254_/B _8178_/B vssd1 vssd1 vccd1 vccd1 _8179_/B sky130_fd_sc_hd__nor2_1
XFILLER_78_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7129_ _6825_/A _6714_/A _7134_/B _7128_/B _7128_/A vssd1 vssd1 vccd1 vccd1 _7131_/A
+ sky130_fd_sc_hd__o32a_1
XFILLER_86_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4830_ _4926_/B vssd1 vssd1 vccd1 vccd1 _4925_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_33_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4761_ _4761_/A vssd1 vssd1 vccd1 vccd1 _8661_/D sky130_fd_sc_hd__clkbuf_1
X_7480_ _7480_/A _7480_/B vssd1 vssd1 vccd1 vccd1 _7481_/B sky130_fd_sc_hd__xnor2_1
X_6500_ _6500_/A vssd1 vssd1 vccd1 vccd1 _8736_/D sky130_fd_sc_hd__clkbuf_1
X_4692_ _7943_/B _8670_/Q _4692_/C _4947_/A vssd1 vssd1 vccd1 vccd1 _4771_/A sky130_fd_sc_hd__or4_2
X_6431_ _6420_/B _6431_/B vssd1 vssd1 vccd1 vccd1 _6431_/X sky130_fd_sc_hd__and2b_1
X_6362_ _6359_/Y _6360_/X _6361_/X vssd1 vssd1 vccd1 vccd1 _6375_/C sky130_fd_sc_hd__o21ai_1
X_8101_ _8214_/A _8100_/X vssd1 vssd1 vccd1 vccd1 _8189_/A sky130_fd_sc_hd__or2b_1
X_5313_ _8674_/Q _5313_/B vssd1 vssd1 vccd1 vccd1 _5313_/X sky130_fd_sc_hd__or2_1
X_6293_ _6293_/A _6293_/B vssd1 vssd1 vccd1 vccd1 _6296_/A sky130_fd_sc_hd__nor2_1
XFILLER_88_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8032_ _8113_/A _8113_/B vssd1 vssd1 vccd1 vccd1 _8114_/A sky130_fd_sc_hd__xnor2_1
X_5244_ _4819_/X _5213_/X _5224_/X _5243_/X _4977_/Y vssd1 vssd1 vccd1 vccd1 _5244_/X
+ sky130_fd_sc_hd__a311o_1
X_5175_ _4964_/X _5171_/X _5174_/X _5164_/X vssd1 vssd1 vccd1 vccd1 _5175_/X sky130_fd_sc_hd__o22a_1
XFILLER_68_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8934_ _8934_/A _4422_/Y vssd1 vssd1 vccd1 vccd1 io_out[21] sky130_fd_sc_hd__ebufn_8
X_7816_ _7745_/A _7902_/B _7828_/B _7904_/A _8155_/A vssd1 vssd1 vccd1 vccd1 _7816_/X
+ sky130_fd_sc_hd__a32o_1
X_7747_ _7754_/A vssd1 vssd1 vccd1 vccd1 _7913_/A sky130_fd_sc_hd__clkbuf_2
X_4959_ _5168_/A _5266_/A vssd1 vssd1 vccd1 vccd1 _4960_/B sky130_fd_sc_hd__nor2_1
X_7678_ _8770_/Q _8667_/Q vssd1 vssd1 vccd1 vccd1 _7678_/X sky130_fd_sc_hd__and2b_1
XFILLER_20_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6629_ _6629_/A _6629_/B vssd1 vssd1 vccd1 vccd1 _6632_/A sky130_fd_sc_hd__nor2_2
XFILLER_10_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6980_ _6980_/A _6980_/B vssd1 vssd1 vccd1 vccd1 _7070_/B sky130_fd_sc_hd__xnor2_1
XFILLER_38_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5931_ _6230_/A vssd1 vssd1 vccd1 vccd1 _6016_/A sky130_fd_sc_hd__clkinv_2
XFILLER_80_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5862_ _5862_/A _5862_/B vssd1 vssd1 vccd1 vccd1 _5937_/B sky130_fd_sc_hd__xnor2_1
X_8650_ _8723_/CLK _8650_/D vssd1 vssd1 vccd1 vccd1 _8650_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5793_ _5792_/A _5792_/B _5792_/C vssd1 vssd1 vccd1 vccd1 _5793_/Y sky130_fd_sc_hd__a21oi_1
X_7601_ _7734_/A _8593_/A _8782_/Q vssd1 vssd1 vccd1 vccd1 _7602_/D sky130_fd_sc_hd__o21a_1
X_8581_ _8582_/A _8582_/B vssd1 vssd1 vccd1 vccd1 _8586_/B sky130_fd_sc_hd__or2_1
X_4813_ _4814_/B _4814_/C _4814_/D _4814_/A vssd1 vssd1 vccd1 vccd1 _4813_/X sky130_fd_sc_hd__a31o_1
X_4744_ _4744_/A _4818_/B vssd1 vssd1 vccd1 vccd1 _5247_/B sky130_fd_sc_hd__nand2_1
X_7532_ _7525_/A _7528_/B _7525_/C _7068_/A vssd1 vssd1 vccd1 vccd1 _7533_/B sky130_fd_sc_hd__a31o_1
X_4675_ _8649_/Q _4674_/B _4640_/X vssd1 vssd1 vccd1 vccd1 _4676_/B sky130_fd_sc_hd__o21ai_1
X_7463_ _7387_/B _7463_/B vssd1 vssd1 vccd1 vccd1 _7463_/X sky130_fd_sc_hd__and2b_1
X_6414_ _5573_/Y _6415_/B _6413_/Y vssd1 vssd1 vccd1 vccd1 _6416_/A sky130_fd_sc_hd__o21a_1
X_7394_ _7451_/A _7394_/B vssd1 vssd1 vccd1 vccd1 _7395_/B sky130_fd_sc_hd__xnor2_2
X_6345_ _6283_/B _6346_/A vssd1 vssd1 vccd1 vccd1 _6345_/X sky130_fd_sc_hd__and2b_1
X_6276_ _6276_/A _6276_/B vssd1 vssd1 vccd1 vccd1 _6280_/A sky130_fd_sc_hd__xor2_2
X_8015_ _8060_/A _8014_/B _8014_/C vssd1 vssd1 vccd1 vccd1 _8016_/C sky130_fd_sc_hd__a21o_1
X_5227_ _5227_/A _5227_/B vssd1 vssd1 vccd1 vccd1 _5235_/A sky130_fd_sc_hd__nor2_2
X_8862__79 vssd1 vssd1 vccd1 vccd1 _8862__79/HI _8971_/A sky130_fd_sc_hd__conb_1
X_5158_ _4701_/A _5154_/X _5156_/X _5197_/D _5157_/X vssd1 vssd1 vccd1 vccd1 _5158_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_84_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5089_ _5188_/B _5163_/A _5157_/B _5226_/A _5066_/A vssd1 vssd1 vccd1 vccd1 _5089_/X
+ sky130_fd_sc_hd__o41a_1
X_8917_ _8917_/A _4400_/Y vssd1 vssd1 vccd1 vccd1 io_out[4] sky130_fd_sc_hd__ebufn_8
XFILLER_37_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8779_ _8783_/CLK _8779_/D vssd1 vssd1 vccd1 vccd1 _8779_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4460_ _4462_/A vssd1 vssd1 vccd1 vccd1 _4460_/Y sky130_fd_sc_hd__inv_2
X_4391_ _4394_/A vssd1 vssd1 vccd1 vccd1 _4391_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6130_ _6132_/A _6132_/B vssd1 vssd1 vccd1 vccd1 _6367_/A sky130_fd_sc_hd__xnor2_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6061_ _6252_/A _6062_/B vssd1 vssd1 vccd1 vccd1 _6178_/A sky130_fd_sc_hd__nor2_1
XFILLER_58_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5012_ _5098_/B _5184_/B _5188_/C _5012_/D vssd1 vssd1 vccd1 vccd1 _5012_/X sky130_fd_sc_hd__or4_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6963_ _6963_/A _6963_/B vssd1 vssd1 vccd1 vccd1 _6967_/B sky130_fd_sc_hd__nor2_1
X_5914_ _5769_/Y _5652_/B _5682_/B _5770_/Y vssd1 vssd1 vccd1 vccd1 _6169_/B sky130_fd_sc_hd__a211o_2
X_6894_ _6894_/A _6894_/B vssd1 vssd1 vccd1 vccd1 _6894_/X sky130_fd_sc_hd__or2_1
X_8702_ _8732_/CLK _8702_/D vssd1 vssd1 vccd1 vccd1 _8702_/Q sky130_fd_sc_hd__dfxtp_1
X_5845_ _5845_/A _5887_/A _5845_/C vssd1 vssd1 vccd1 vccd1 _5887_/B sky130_fd_sc_hd__nand3_1
XFILLER_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8633_ _8732_/CLK _8633_/D vssd1 vssd1 vccd1 vccd1 _8633_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5776_ _6107_/A _5916_/B _6107_/B vssd1 vssd1 vccd1 vccd1 _5777_/B sky130_fd_sc_hd__a21oi_1
X_8564_ _8554_/X _8555_/Y _8558_/X _8561_/Y _8563_/Y vssd1 vssd1 vccd1 vccd1 _8565_/D
+ sky130_fd_sc_hd__a2111o_1
X_8495_ _8422_/A _8422_/B _8494_/X vssd1 vssd1 vccd1 vccd1 _8500_/A sky130_fd_sc_hd__a21o_1
X_4727_ _4733_/B _4733_/C vssd1 vssd1 vccd1 vccd1 _4734_/B sky130_fd_sc_hd__and2_1
X_7515_ _7515_/A _7515_/B _7518_/A vssd1 vssd1 vccd1 vccd1 _7516_/B sky130_fd_sc_hd__and3_1
X_4658_ _4661_/C _4658_/B vssd1 vssd1 vccd1 vccd1 _8643_/D sky130_fd_sc_hd__nor2_1
X_7446_ _7446_/A _7396_/A vssd1 vssd1 vccd1 vccd1 _7446_/X sky130_fd_sc_hd__or2b_1
XFILLER_103_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4589_ _8682_/Q _4595_/B vssd1 vssd1 vccd1 vccd1 _4590_/A sky130_fd_sc_hd__and2_1
XFILLER_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7377_ _7377_/A vssd1 vssd1 vccd1 vccd1 _7388_/S sky130_fd_sc_hd__clkbuf_2
X_6328_ _5634_/A _5634_/C _5735_/X vssd1 vssd1 vccd1 vccd1 _6330_/A sky130_fd_sc_hd__a21o_1
XFILLER_103_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6259_ _6259_/A _6259_/B vssd1 vssd1 vccd1 vccd1 _6268_/A sky130_fd_sc_hd__and2_1
XFILLER_67_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5630_ _5630_/A vssd1 vssd1 vccd1 vccd1 _6092_/A sky130_fd_sc_hd__clkbuf_2
X_5561_ _5615_/A _5561_/B vssd1 vssd1 vccd1 vccd1 _5608_/A sky130_fd_sc_hd__nor2_4
X_8280_ _8280_/A _8280_/B _8280_/C _8280_/D vssd1 vssd1 vccd1 vccd1 _8282_/A sky130_fd_sc_hd__and4_1
X_5492_ _6621_/B _8707_/Q vssd1 vssd1 vccd1 vccd1 _5493_/A sky130_fd_sc_hd__or2b_1
X_7300_ _7300_/A vssd1 vssd1 vccd1 vccd1 _7309_/B sky130_fd_sc_hd__clkbuf_2
X_4512_ _4877_/B vssd1 vssd1 vccd1 vccd1 _4778_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7231_ _7231_/A _7231_/B vssd1 vssd1 vccd1 vccd1 _7327_/B sky130_fd_sc_hd__xnor2_1
X_4443_ _4444_/A vssd1 vssd1 vccd1 vccd1 _4443_/Y sky130_fd_sc_hd__inv_2
X_4374_ _4376_/A vssd1 vssd1 vccd1 vccd1 _4374_/Y sky130_fd_sc_hd__inv_2
X_7162_ _7062_/A _7062_/B _7161_/X vssd1 vssd1 vccd1 vccd1 _7243_/A sky130_fd_sc_hd__a21bo_1
X_6113_ _6157_/A _6113_/B vssd1 vssd1 vccd1 vccd1 _6116_/A sky130_fd_sc_hd__xor2_1
X_7093_ _7093_/A _7093_/B vssd1 vssd1 vccd1 vccd1 _7097_/B sky130_fd_sc_hd__xor2_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6044_ _6044_/A _6044_/B vssd1 vssd1 vccd1 vccd1 _6045_/B sky130_fd_sc_hd__xor2_2
X_8832__49 vssd1 vssd1 vccd1 vccd1 _8832__49/HI _8941_/A sky130_fd_sc_hd__conb_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7995_ _8063_/B _7994_/C _7994_/A vssd1 vssd1 vccd1 vccd1 _8002_/B sky130_fd_sc_hd__a21o_1
XFILLER_54_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6946_ _7416_/A _7050_/A vssd1 vssd1 vccd1 vccd1 _6947_/B sky130_fd_sc_hd__nand2_1
XFILLER_26_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6877_ _6877_/A _6877_/B vssd1 vssd1 vccd1 vccd1 _6922_/B sky130_fd_sc_hd__xor2_2
X_5828_ _6263_/A _5980_/A _5827_/X vssd1 vssd1 vccd1 vccd1 _5829_/B sky130_fd_sc_hd__a21oi_1
X_8616_ _8615_/A _8615_/C _8615_/B vssd1 vssd1 vccd1 vccd1 _8616_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_22_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5759_ _5811_/B _5811_/C _5811_/A vssd1 vssd1 vccd1 vccd1 _5760_/D sky130_fd_sc_hd__a21o_1
X_8547_ _8547_/A _8547_/B _8547_/C vssd1 vssd1 vccd1 vccd1 _8565_/B sky130_fd_sc_hd__and3_1
X_8478_ _8491_/A _8478_/B vssd1 vssd1 vccd1 vccd1 _8479_/B sky130_fd_sc_hd__and2_1
X_7429_ _7505_/A _7505_/B vssd1 vssd1 vccd1 vccd1 _7430_/B sky130_fd_sc_hd__xor2_2
XFILLER_89_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6800_ _6801_/A _6801_/B _6801_/C vssd1 vssd1 vccd1 vccd1 _6802_/A sky130_fd_sc_hd__a21o_1
X_7780_ _8349_/A vssd1 vssd1 vccd1 vccd1 _8348_/A sky130_fd_sc_hd__clkbuf_2
X_4992_ _5168_/A vssd1 vssd1 vccd1 vccd1 _5176_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_51_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6731_ _6970_/A _6970_/B vssd1 vssd1 vccd1 vccd1 _6891_/A sky130_fd_sc_hd__or2b_1
XFILLER_31_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6662_ _8764_/Q _7794_/B vssd1 vssd1 vccd1 vccd1 _6662_/X sky130_fd_sc_hd__and2b_1
X_8401_ _8434_/A _8401_/B vssd1 vssd1 vccd1 vccd1 _8411_/B sky130_fd_sc_hd__xnor2_2
X_5613_ _5688_/A vssd1 vssd1 vccd1 vccd1 _5727_/A sky130_fd_sc_hd__inv_2
X_8332_ _8198_/A _8417_/A _8332_/C vssd1 vssd1 vccd1 vccd1 _8417_/B sky130_fd_sc_hd__nand3b_1
X_6593_ _6593_/A _7576_/B _7583_/B vssd1 vssd1 vccd1 vccd1 _6593_/X sky130_fd_sc_hd__and3_1
X_5544_ _5544_/A _5544_/B vssd1 vssd1 vccd1 vccd1 _5554_/B sky130_fd_sc_hd__and2_2
X_8263_ _8382_/A _8263_/B vssd1 vssd1 vccd1 vccd1 _8386_/A sky130_fd_sc_hd__nand2_1
X_5475_ _5480_/A _5475_/B _5475_/C vssd1 vssd1 vccd1 vccd1 _5485_/S sky130_fd_sc_hd__nand3_2
X_4426_ _4426_/A vssd1 vssd1 vccd1 vccd1 _4431_/A sky130_fd_sc_hd__buf_8
X_8194_ _8236_/C _8194_/B vssd1 vssd1 vccd1 vccd1 _8197_/A sky130_fd_sc_hd__xnor2_1
X_7214_ _7214_/A _7214_/B vssd1 vssd1 vccd1 vccd1 _7215_/B sky130_fd_sc_hd__xnor2_1
X_7145_ _7151_/A _7145_/B vssd1 vssd1 vccd1 vccd1 _7146_/A sky130_fd_sc_hd__nor2_1
XFILLER_98_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4357_ _4481_/A vssd1 vssd1 vccd1 vccd1 _4489_/A sky130_fd_sc_hd__buf_6
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7076_ _7100_/A _7083_/B vssd1 vssd1 vccd1 vccd1 _7098_/A sky130_fd_sc_hd__xor2_1
XFILLER_104_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6027_ _6027_/A _6027_/B vssd1 vssd1 vccd1 vccd1 _6028_/B sky130_fd_sc_hd__nor2_1
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7978_ _8138_/A _8139_/A vssd1 vssd1 vccd1 vccd1 _7979_/B sky130_fd_sc_hd__nand2_1
XFILLER_14_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6929_ _7019_/A _6928_/X _6873_/B vssd1 vssd1 vccd1 vccd1 _7028_/A sky130_fd_sc_hd__a21oi_2
XFILLER_42_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_49_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5260_ _5258_/X _5259_/X _4974_/X vssd1 vssd1 vccd1 vccd1 _5296_/C sky130_fd_sc_hd__o21a_1
XFILLER_102_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5191_ _5274_/A _5127_/A _5188_/X _5190_/X vssd1 vssd1 vccd1 vccd1 _5192_/D sky130_fd_sc_hd__o31a_1
XFILLER_95_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8802__19 vssd1 vssd1 vccd1 vccd1 _8802__19/HI _8897_/A sky130_fd_sc_hd__conb_1
XFILLER_68_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8950_ _8950_/A _4444_/Y vssd1 vssd1 vccd1 vccd1 io_out[37] sky130_fd_sc_hd__ebufn_8
XFILLER_83_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7901_ _7924_/A _8158_/A _7802_/B _7907_/B vssd1 vssd1 vccd1 vccd1 _7910_/A sky130_fd_sc_hd__a31o_1
XFILLER_36_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8881_ _8881_/A _4489_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[0] sky130_fd_sc_hd__ebufn_8
X_7832_ _7998_/A _8163_/A vssd1 vssd1 vccd1 vccd1 _7833_/C sky130_fd_sc_hd__nand2_1
XFILLER_34_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7763_ _8024_/A _8092_/A vssd1 vssd1 vccd1 vccd1 _8332_/C sky130_fd_sc_hd__or2_1
XFILLER_24_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4975_ _4819_/X _4962_/X _4972_/X _4974_/X vssd1 vssd1 vccd1 vccd1 _4975_/X sky130_fd_sc_hd__o211a_1
XFILLER_11_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6714_ _6714_/A _6714_/B vssd1 vssd1 vccd1 vccd1 _7078_/B sky130_fd_sc_hd__xor2_2
X_7694_ _8330_/A vssd1 vssd1 vccd1 vccd1 _8325_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6645_ _6645_/A _6645_/B vssd1 vssd1 vccd1 vccd1 _6646_/A sky130_fd_sc_hd__nand2_1
X_6576_ _8750_/Q vssd1 vssd1 vccd1 vccd1 _6577_/A sky130_fd_sc_hd__inv_2
X_5527_ _5527_/A vssd1 vssd1 vccd1 vccd1 _6107_/A sky130_fd_sc_hd__clkbuf_2
X_8315_ _8315_/A _8315_/B vssd1 vssd1 vccd1 vccd1 _8554_/B sky130_fd_sc_hd__nor2_1
X_8246_ _8180_/A _8246_/B vssd1 vssd1 vccd1 vccd1 _8246_/X sky130_fd_sc_hd__and2b_1
XFILLER_59_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5458_ _5458_/A _5458_/B vssd1 vssd1 vccd1 vccd1 _5460_/A sky130_fd_sc_hd__nor2_1
X_4409_ _4413_/A vssd1 vssd1 vccd1 vccd1 _4409_/Y sky130_fd_sc_hd__inv_2
X_8177_ _8177_/A _8177_/B vssd1 vssd1 vccd1 vccd1 _8178_/B sky130_fd_sc_hd__nor2_1
X_5389_ _5395_/C _5389_/B _5389_/C vssd1 vssd1 vccd1 vccd1 _5390_/A sky130_fd_sc_hd__and3b_1
XFILLER_86_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7128_ _7128_/A _7128_/B vssd1 vssd1 vccd1 vccd1 _7134_/B sky130_fd_sc_hd__xnor2_1
XFILLER_101_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7059_ _7163_/B _7059_/B vssd1 vssd1 vccd1 vccd1 _7060_/B sky130_fd_sc_hd__xnor2_1
XFILLER_46_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8789__6 vssd1 vssd1 vccd1 vccd1 _8789__6/HI _8884_/A sky130_fd_sc_hd__conb_1
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8868__85 vssd1 vssd1 vccd1 vccd1 _8868__85/HI _8977_/A sky130_fd_sc_hd__conb_1
XFILLER_40_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4760_ _4760_/A _4760_/B _4760_/C vssd1 vssd1 vccd1 vccd1 _4761_/A sky130_fd_sc_hd__and3_1
XFILLER_14_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4691_ _4872_/B _4762_/A _4812_/B vssd1 vssd1 vccd1 vccd1 _4947_/A sky130_fd_sc_hd__or3_4
X_6430_ _5450_/X _6429_/Y _6427_/A _4616_/B vssd1 vssd1 vccd1 vccd1 _8723_/D sky130_fd_sc_hd__o2bb2a_1
X_6361_ _6361_/A _6361_/B vssd1 vssd1 vccd1 vccd1 _6361_/X sky130_fd_sc_hd__xor2_1
X_8100_ _8099_/A _8327_/A _8099_/D _8099_/C vssd1 vssd1 vccd1 vccd1 _8100_/X sky130_fd_sc_hd__a31o_1
X_5312_ _8715_/Q _5307_/X _5310_/X _5311_/X vssd1 vssd1 vccd1 vccd1 _8673_/D sky130_fd_sc_hd__o211a_1
X_6292_ _6292_/A _6292_/B vssd1 vssd1 vccd1 vccd1 _6361_/B sky130_fd_sc_hd__xor2_1
X_8031_ _8111_/A _8031_/B vssd1 vssd1 vccd1 vccd1 _8113_/B sky130_fd_sc_hd__nor2_1
X_5243_ _5224_/C _5242_/X _5170_/A vssd1 vssd1 vccd1 vccd1 _5243_/X sky130_fd_sc_hd__o21a_1
X_5174_ _5174_/A _5174_/B _5174_/C vssd1 vssd1 vccd1 vccd1 _5174_/X sky130_fd_sc_hd__or3_1
XFILLER_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8933_ _8933_/A _4421_/Y vssd1 vssd1 vccd1 vccd1 io_out[20] sky130_fd_sc_hd__ebufn_8
XFILLER_101_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7815_ _8155_/C vssd1 vssd1 vccd1 vccd1 _7828_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_52_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7746_ _7788_/A _7788_/B vssd1 vssd1 vccd1 vccd1 _7754_/A sky130_fd_sc_hd__xnor2_2
X_4958_ _5210_/A vssd1 vssd1 vccd1 vccd1 _5168_/A sky130_fd_sc_hd__clkbuf_2
X_7677_ _7762_/A _7708_/B _7676_/X vssd1 vssd1 vccd1 vccd1 _7681_/A sky130_fd_sc_hd__a21o_1
X_4889_ _4935_/A _4889_/B vssd1 vssd1 vccd1 vccd1 _5156_/A sky130_fd_sc_hd__nor2_1
XFILLER_20_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6628_ _6627_/B _6628_/B vssd1 vssd1 vccd1 vccd1 _6629_/B sky130_fd_sc_hd__and2b_1
X_6559_ _6758_/A _6557_/X _6590_/A _8754_/Q vssd1 vssd1 vccd1 vccd1 _6560_/B sky130_fd_sc_hd__a31oi_1
XFILLER_79_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8229_ _8229_/A _8229_/B vssd1 vssd1 vccd1 vccd1 _8229_/Y sky130_fd_sc_hd__nor2_1
XFILLER_10_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5930_ _5943_/B _5946_/B vssd1 vssd1 vccd1 vccd1 _5933_/A sky130_fd_sc_hd__or2b_1
XFILLER_53_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5861_ _5922_/A _5861_/B vssd1 vssd1 vccd1 vccd1 _5862_/B sky130_fd_sc_hd__nor2_1
X_7600_ _8785_/Q vssd1 vssd1 vccd1 vccd1 _7602_/A sky130_fd_sc_hd__clkbuf_2
X_5792_ _5792_/A _5792_/B _5792_/C vssd1 vssd1 vccd1 vccd1 _5792_/X sky130_fd_sc_hd__and3_1
X_8580_ _6387_/X _8573_/X _8578_/X _8579_/Y vssd1 vssd1 vccd1 vccd1 _8776_/D sky130_fd_sc_hd__a31oi_1
X_4812_ _4877_/C _4812_/B vssd1 vssd1 vccd1 vccd1 _4814_/D sky130_fd_sc_hd__nor2_1
X_4743_ _4740_/A _4742_/A _4742_/Y _4705_/X vssd1 vssd1 vccd1 vccd1 _8657_/D sky130_fd_sc_hd__o211a_1
X_7531_ _7525_/X _7526_/Y _7529_/Y _7530_/Y vssd1 vssd1 vccd1 vccd1 _7540_/B sky130_fd_sc_hd__o211ai_4
X_7462_ _7462_/A _7462_/B vssd1 vssd1 vccd1 vccd1 _7465_/B sky130_fd_sc_hd__nand2_1
X_4674_ _8649_/Q _4674_/B vssd1 vssd1 vccd1 vccd1 _4678_/B sky130_fd_sc_hd__and2_1
X_6413_ _6413_/A _6413_/B vssd1 vssd1 vccd1 vccd1 _6413_/Y sky130_fd_sc_hd__nand2_1
X_7393_ _7228_/A _7391_/Y _7450_/S vssd1 vssd1 vccd1 vccd1 _7394_/B sky130_fd_sc_hd__mux2_1
X_6344_ _6242_/A _6342_/Y _6343_/X vssd1 vssd1 vccd1 vccd1 _6348_/A sky130_fd_sc_hd__a21o_1
XFILLER_88_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6275_ _5827_/X _6274_/Y _6275_/S vssd1 vssd1 vccd1 vccd1 _6276_/B sky130_fd_sc_hd__mux2_1
XFILLER_88_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8014_ _8060_/A _8014_/B _8014_/C vssd1 vssd1 vccd1 vccd1 _8060_/B sky130_fd_sc_hd__nand3_1
X_5226_ _5226_/A _5227_/B vssd1 vssd1 vccd1 vccd1 _5226_/Y sky130_fd_sc_hd__nor2_1
XFILLER_102_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5157_ _5157_/A _5157_/B _5251_/B _5157_/D vssd1 vssd1 vccd1 vccd1 _5157_/X sky130_fd_sc_hd__or4_1
XFILLER_96_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5088_ _5088_/A _5088_/B vssd1 vssd1 vccd1 vccd1 _5226_/A sky130_fd_sc_hd__nand2_1
XFILLER_29_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8916_ _8916_/A _4399_/Y vssd1 vssd1 vccd1 vccd1 io_out[3] sky130_fd_sc_hd__ebufn_8
XFILLER_56_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8778_ _8778_/CLK _8778_/D vssd1 vssd1 vccd1 vccd1 _8778_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7729_ _8780_/Q _7729_/B vssd1 vssd1 vccd1 vccd1 _7729_/X sky130_fd_sc_hd__and2b_1
XFILLER_4_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8838__55 vssd1 vssd1 vccd1 vccd1 _8838__55/HI _8947_/A sky130_fd_sc_hd__conb_1
XFILLER_97_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4390_ _4394_/A vssd1 vssd1 vccd1 vccd1 _4390_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6060_ _6249_/A _6059_/X _6014_/Y vssd1 vssd1 vccd1 vccd1 _6062_/B sky130_fd_sc_hd__a21o_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5011_ _5283_/A _5157_/A _5283_/C _5172_/C vssd1 vssd1 vccd1 vccd1 _5012_/D sky130_fd_sc_hd__or4_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6962_ _6786_/A _7119_/A _6767_/C vssd1 vssd1 vccd1 vccd1 _6963_/B sky130_fd_sc_hd__a21oi_1
X_5913_ _5913_/A _5925_/B vssd1 vssd1 vccd1 vccd1 _6144_/A sky130_fd_sc_hd__nand2_1
X_6893_ _6982_/A _6982_/B _6892_/Y vssd1 vssd1 vccd1 vccd1 _6955_/A sky130_fd_sc_hd__a21oi_1
X_8701_ _8732_/CLK _8701_/D vssd1 vssd1 vccd1 vccd1 _8701_/Q sky130_fd_sc_hd__dfxtp_1
X_5844_ _5888_/B _5843_/C _5843_/A vssd1 vssd1 vccd1 vccd1 _5845_/C sky130_fd_sc_hd__a21o_1
XFILLER_22_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8632_ _8730_/CLK _8632_/D vssd1 vssd1 vccd1 vccd1 _8632_/Q sky130_fd_sc_hd__dfxtp_1
X_8563_ _8563_/A _8563_/B vssd1 vssd1 vccd1 vccd1 _8563_/Y sky130_fd_sc_hd__nor2_1
X_5775_ _5775_/A vssd1 vssd1 vccd1 vccd1 _6107_/B sky130_fd_sc_hd__buf_2
X_7514_ _7514_/A _7514_/B vssd1 vssd1 vccd1 vccd1 _7552_/A sky130_fd_sc_hd__xnor2_4
XFILLER_21_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8494_ _8421_/A _8494_/B vssd1 vssd1 vccd1 vccd1 _8494_/X sky130_fd_sc_hd__and2b_1
X_4726_ _4733_/B _4733_/C vssd1 vssd1 vccd1 vccd1 _4818_/A sky130_fd_sc_hd__nor2_1
X_4657_ _8643_/Q _4656_/B _4640_/X vssd1 vssd1 vccd1 vccd1 _4658_/B sky130_fd_sc_hd__o21ai_1
X_7445_ _7374_/A _7374_/B _7444_/X vssd1 vssd1 vccd1 vccd1 _7456_/A sky130_fd_sc_hd__a21oi_1
X_7376_ _7272_/A _7409_/B _7272_/C _7278_/A vssd1 vssd1 vccd1 vccd1 _7396_/A sky130_fd_sc_hd__a31o_1
X_4588_ _4588_/A vssd1 vssd1 vccd1 vccd1 _8935_/A sky130_fd_sc_hd__clkbuf_1
X_6327_ _6281_/A _6281_/B _6326_/Y vssd1 vssd1 vccd1 vccd1 _6331_/A sky130_fd_sc_hd__a21oi_1
XFILLER_1_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6258_ _6209_/A _6209_/B _6208_/A vssd1 vssd1 vccd1 vccd1 _6346_/A sky130_fd_sc_hd__a21oi_1
XFILLER_88_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6189_ _6248_/A _6189_/B vssd1 vssd1 vccd1 vccd1 _6209_/A sky130_fd_sc_hd__xnor2_1
XFILLER_57_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5209_ _5209_/A _5209_/B vssd1 vssd1 vccd1 vccd1 _5210_/B sky130_fd_sc_hd__nor2_1
XFILLER_57_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5560_ _6655_/B _8722_/Q vssd1 vssd1 vccd1 vccd1 _5561_/B sky130_fd_sc_hd__and2b_1
X_5491_ _7656_/B vssd1 vssd1 vccd1 vccd1 _5491_/X sky130_fd_sc_hd__buf_2
X_4511_ _4878_/B vssd1 vssd1 vccd1 vccd1 _4877_/B sky130_fd_sc_hd__clkbuf_1
X_7230_ _7230_/A _7230_/B vssd1 vssd1 vccd1 vccd1 _7231_/B sky130_fd_sc_hd__xnor2_1
XFILLER_7_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4442_ _4444_/A vssd1 vssd1 vccd1 vccd1 _4442_/Y sky130_fd_sc_hd__inv_2
X_4373_ _4376_/A vssd1 vssd1 vccd1 vccd1 _4373_/Y sky130_fd_sc_hd__inv_2
X_7161_ _7161_/A _7063_/A vssd1 vssd1 vccd1 vccd1 _7161_/X sky130_fd_sc_hd__or2b_1
X_6112_ _6156_/A _6156_/B vssd1 vssd1 vccd1 vccd1 _6113_/B sky130_fd_sc_hd__xor2_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7092_ _7092_/A _7092_/B vssd1 vssd1 vccd1 vccd1 _7093_/A sky130_fd_sc_hd__nand2_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6043_ _6043_/A _6043_/B vssd1 vssd1 vccd1 vccd1 _6044_/B sky130_fd_sc_hd__nand2_1
XFILLER_85_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7994_ _7994_/A _8063_/B _7994_/C vssd1 vssd1 vccd1 vccd1 _8061_/A sky130_fd_sc_hd__nand3_1
XFILLER_81_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6945_ _7212_/A vssd1 vssd1 vccd1 vccd1 _7373_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_26_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_2_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
X_6876_ _6876_/A _6862_/X vssd1 vssd1 vccd1 vccd1 _6877_/B sky130_fd_sc_hd__or2b_1
X_5827_ _5827_/A vssd1 vssd1 vccd1 vccd1 _5827_/X sky130_fd_sc_hd__clkbuf_2
X_8615_ _8615_/A _8615_/B _8615_/C vssd1 vssd1 vccd1 vccd1 _8627_/S sky130_fd_sc_hd__or3_1
X_5758_ _5811_/A _5811_/B _5811_/C vssd1 vssd1 vccd1 vccd1 _5760_/C sky130_fd_sc_hd__nand3_1
X_8546_ _8547_/A _8547_/B _8547_/C vssd1 vssd1 vccd1 vccd1 _8565_/A sky130_fd_sc_hd__a21oi_1
X_8477_ _8477_/A _8477_/B _8477_/C vssd1 vssd1 vccd1 vccd1 _8478_/B sky130_fd_sc_hd__or3_1
XFILLER_5_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4709_ _5221_/A vssd1 vssd1 vccd1 vccd1 _4946_/A sky130_fd_sc_hd__clkbuf_2
X_5689_ _5991_/A _5701_/B vssd1 vssd1 vccd1 vccd1 _5702_/A sky130_fd_sc_hd__nor2_1
X_7428_ _7321_/A _7321_/B _7427_/Y vssd1 vssd1 vccd1 vccd1 _7505_/B sky130_fd_sc_hd__o21ai_2
X_8808__25 vssd1 vssd1 vccd1 vccd1 _8808__25/HI _8903_/A sky130_fd_sc_hd__conb_1
X_7359_ _7366_/A vssd1 vssd1 vccd1 vccd1 _7508_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_1_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6730_ _6723_/X _6728_/Y _6729_/X vssd1 vssd1 vccd1 vccd1 _6970_/B sky130_fd_sc_hd__o21a_1
X_4991_ _5136_/A _4894_/B _4946_/A vssd1 vssd1 vccd1 vccd1 _4991_/Y sky130_fd_sc_hd__o21ai_1
X_6661_ _6670_/A _6670_/B _6703_/B _6617_/A vssd1 vssd1 vccd1 vccd1 _6695_/B sky130_fd_sc_hd__a211o_1
X_8400_ _8435_/A _8435_/B vssd1 vssd1 vccd1 vccd1 _8401_/B sky130_fd_sc_hd__xor2_2
X_5612_ _6262_/A _5720_/B vssd1 vssd1 vccd1 vccd1 _5627_/A sky130_fd_sc_hd__xnor2_1
X_6592_ _7587_/B vssd1 vssd1 vccd1 vccd1 _7583_/B sky130_fd_sc_hd__clkbuf_2
X_8331_ _8332_/C _8417_/A _7839_/B vssd1 vssd1 vccd1 vccd1 _8333_/B sky130_fd_sc_hd__a21o_1
X_5543_ _5505_/A _5505_/B _5508_/X _5518_/X _5509_/A vssd1 vssd1 vccd1 vccd1 _5544_/B
+ sky130_fd_sc_hd__a311o_1
X_8262_ _8262_/A _8263_/B vssd1 vssd1 vccd1 vccd1 _8264_/B sky130_fd_sc_hd__or2_1
X_5474_ _5480_/A _5475_/B _5475_/C vssd1 vssd1 vccd1 vccd1 _5474_/X sky130_fd_sc_hd__a21o_1
X_4425_ _4425_/A vssd1 vssd1 vccd1 vccd1 _4425_/Y sky130_fd_sc_hd__inv_2
X_8193_ _8239_/A _8418_/A _8192_/Y vssd1 vssd1 vccd1 vccd1 _8194_/B sky130_fd_sc_hd__o21bai_2
X_7213_ _7334_/A _7213_/B vssd1 vssd1 vccd1 vccd1 _7214_/B sky130_fd_sc_hd__and2_1
X_4356_ input1/X vssd1 vssd1 vccd1 vccd1 _4481_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7144_ _7151_/A _7145_/B _7146_/B vssd1 vssd1 vccd1 vccd1 _7515_/B sky130_fd_sc_hd__or3_1
XFILLER_98_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7075_ _7075_/A _7075_/B vssd1 vssd1 vccd1 vccd1 _7083_/B sky130_fd_sc_hd__xor2_1
X_6026_ _6027_/A _6027_/B vssd1 vssd1 vccd1 vccd1 _6119_/B sky130_fd_sc_hd__and2_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7977_ _8053_/A _7977_/B vssd1 vssd1 vccd1 vccd1 _8139_/B sky130_fd_sc_hd__or2_1
XFILLER_27_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6928_ _6765_/A _6836_/A _6792_/B _6863_/C _7020_/A vssd1 vssd1 vccd1 vccd1 _6928_/X
+ sky130_fd_sc_hd__a32o_1
X_6859_ _7378_/A vssd1 vssd1 vccd1 vccd1 _7489_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_50_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8529_ _8456_/A _8456_/B _8528_/Y vssd1 vssd1 vccd1 vccd1 _8532_/A sky130_fd_sc_hd__o21a_1
XFILLER_6_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8799__16 vssd1 vssd1 vccd1 vccd1 _8799__16/HI _8894_/A sky130_fd_sc_hd__conb_1
XFILLER_68_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5190_ _5190_/A _5274_/A _5190_/C _5190_/D vssd1 vssd1 vccd1 vccd1 _5190_/X sky130_fd_sc_hd__or4_1
XFILLER_95_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7900_ _8155_/A _7904_/A _7996_/A vssd1 vssd1 vccd1 vccd1 _7907_/B sky130_fd_sc_hd__and3_1
XFILLER_55_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7831_ _7831_/A _7831_/B vssd1 vssd1 vccd1 vccd1 _7834_/A sky130_fd_sc_hd__xnor2_1
XFILLER_36_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7762_ _7762_/A _7762_/B vssd1 vssd1 vccd1 vccd1 _7940_/A sky130_fd_sc_hd__nand2_1
X_4974_ _5224_/A vssd1 vssd1 vccd1 vccd1 _4974_/X sky130_fd_sc_hd__clkbuf_2
X_7693_ _7693_/A vssd1 vssd1 vccd1 vccd1 _8330_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6713_ _6713_/A _6713_/B vssd1 vssd1 vccd1 vccd1 _6714_/B sky130_fd_sc_hd__nand2_1
X_6644_ _6644_/A _6644_/B vssd1 vssd1 vccd1 vccd1 _6651_/A sky130_fd_sc_hd__nand2_1
XFILLER_50_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6575_ _6628_/B _6583_/B vssd1 vssd1 vccd1 vccd1 _6578_/A sky130_fd_sc_hd__nor2_1
X_5526_ _5552_/A _5526_/B vssd1 vssd1 vccd1 vccd1 _5527_/A sky130_fd_sc_hd__xor2_2
X_8314_ _8562_/B _8562_/C _8310_/Y _8562_/A vssd1 vssd1 vccd1 vccd1 _8549_/B sky130_fd_sc_hd__a211o_1
X_8245_ _8245_/A _8245_/B vssd1 vssd1 vccd1 vccd1 _8286_/A sky130_fd_sc_hd__xor2_2
X_5457_ _5456_/B _5478_/B vssd1 vssd1 vccd1 vccd1 _5458_/B sky130_fd_sc_hd__and2b_1
X_4408_ _4426_/A vssd1 vssd1 vccd1 vccd1 _4413_/A sky130_fd_sc_hd__buf_4
X_8176_ _8177_/A _8177_/B vssd1 vssd1 vccd1 vccd1 _8254_/B sky130_fd_sc_hd__and2_1
X_5388_ _6528_/C _8694_/Q _5381_/B _8696_/Q vssd1 vssd1 vccd1 vccd1 _5389_/C sky130_fd_sc_hd__a31o_1
XFILLER_86_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7127_ _7127_/A _7127_/B vssd1 vssd1 vccd1 vccd1 _7128_/B sky130_fd_sc_hd__nand2_1
XFILLER_86_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7058_ _7373_/A _7058_/B vssd1 vssd1 vccd1 vccd1 _7059_/B sky130_fd_sc_hd__xnor2_1
XFILLER_101_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6009_ _6009_/A _6009_/B vssd1 vssd1 vccd1 vccd1 _6055_/B sky130_fd_sc_hd__xnor2_2
XFILLER_75_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4690_ _4878_/A _4878_/B vssd1 vssd1 vccd1 vccd1 _4812_/B sky130_fd_sc_hd__nand2_1
X_6360_ _6360_/A _6360_/B _6360_/C vssd1 vssd1 vccd1 vccd1 _6360_/X sky130_fd_sc_hd__and3_1
X_5311_ _5335_/A vssd1 vssd1 vccd1 vccd1 _5311_/X sky130_fd_sc_hd__clkbuf_2
X_6291_ _6304_/A _6291_/B vssd1 vssd1 vccd1 vccd1 _6292_/B sky130_fd_sc_hd__and2_1
X_8030_ _8044_/A _8030_/B _8034_/A vssd1 vssd1 vccd1 vccd1 _8031_/B sky130_fd_sc_hd__nor3_1
X_5242_ _5224_/A _5232_/X _5241_/X vssd1 vssd1 vccd1 vccd1 _5242_/X sky130_fd_sc_hd__o21a_1
X_5173_ _5261_/D _5173_/B vssd1 vssd1 vccd1 vccd1 _5174_/C sky130_fd_sc_hd__or2_1
XFILLER_96_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput1 active vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_6
XFILLER_96_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8932_ _8932_/A _4419_/Y vssd1 vssd1 vccd1 vccd1 io_out[19] sky130_fd_sc_hd__ebufn_8
XFILLER_83_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7814_ _8155_/B vssd1 vssd1 vccd1 vccd1 _7902_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_24_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7745_ _7745_/A vssd1 vssd1 vccd1 vccd1 _7934_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_61_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4957_ _4957_/A vssd1 vssd1 vccd1 vccd1 _5149_/C sky130_fd_sc_hd__clkbuf_2
X_7676_ _8769_/Q _8666_/Q vssd1 vssd1 vccd1 vccd1 _7676_/X sky130_fd_sc_hd__and2b_1
X_4888_ _4889_/B _4910_/B _4887_/X vssd1 vssd1 vccd1 vccd1 _5272_/B sky130_fd_sc_hd__o21ai_4
XFILLER_20_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6627_ _8750_/Q _6627_/B vssd1 vssd1 vccd1 vccd1 _6629_/A sky130_fd_sc_hd__and2b_1
X_6558_ _6593_/A _6588_/B vssd1 vssd1 vccd1 vccd1 _6590_/A sky130_fd_sc_hd__or2_1
X_5509_ _5509_/A _5508_/X vssd1 vssd1 vccd1 vccd1 _5530_/B sky130_fd_sc_hd__nor2b_4
X_6489_ _8733_/Q _6492_/C vssd1 vssd1 vccd1 vccd1 _6491_/A sky130_fd_sc_hd__and2_1
X_8228_ _8228_/A vssd1 vssd1 vccd1 vccd1 _8228_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8159_ _8158_/B _8158_/C _8248_/B vssd1 vssd1 vccd1 vccd1 _8272_/B sky130_fd_sc_hd__a21oi_1
XFILLER_87_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8791__8 vssd1 vssd1 vccd1 vccd1 _8791__8/HI _8886_/A sky130_fd_sc_hd__conb_1
XFILLER_47_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5860_ _5936_/A _5936_/B vssd1 vssd1 vccd1 vccd1 _5937_/A sky130_fd_sc_hd__xnor2_1
X_4811_ _4811_/A vssd1 vssd1 vccd1 vccd1 _8670_/D sky130_fd_sc_hd__clkbuf_1
X_5791_ _5884_/A _5791_/B vssd1 vssd1 vccd1 vccd1 _5792_/C sky130_fd_sc_hd__nor2_1
X_4742_ _4742_/A _5296_/A vssd1 vssd1 vccd1 vccd1 _4742_/Y sky130_fd_sc_hd__nand2_1
X_7530_ _7530_/A _7530_/B vssd1 vssd1 vccd1 vccd1 _7530_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_21_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4673_ _4673_/A vssd1 vssd1 vccd1 vccd1 _8648_/D sky130_fd_sc_hd__clkbuf_1
X_7461_ _7461_/A _7461_/B vssd1 vssd1 vccd1 vccd1 _7465_/A sky130_fd_sc_hd__nand2_1
X_6412_ _6409_/A _5449_/X _5450_/A _6411_/X vssd1 vssd1 vccd1 vccd1 _8720_/D sky130_fd_sc_hd__a22o_1
X_7392_ _7392_/A _7392_/B vssd1 vssd1 vccd1 vccd1 _7450_/S sky130_fd_sc_hd__xor2_1
X_6343_ _6239_/B _6343_/B vssd1 vssd1 vccd1 vccd1 _6343_/X sky130_fd_sc_hd__and2b_1
X_6274_ _6274_/A _6274_/B vssd1 vssd1 vccd1 vccd1 _6274_/Y sky130_fd_sc_hd__nor2_1
XFILLER_88_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8013_ _8083_/A _8013_/B vssd1 vssd1 vccd1 vccd1 _8014_/C sky130_fd_sc_hd__xnor2_1
XFILLER_69_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5225_ _5250_/B _5225_/B _5285_/B _5234_/A vssd1 vssd1 vccd1 vccd1 _5225_/X sky130_fd_sc_hd__or4_1
XFILLER_69_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5156_ _5156_/A _5156_/B _5157_/D vssd1 vssd1 vccd1 vccd1 _5156_/X sky130_fd_sc_hd__or3_1
X_5087_ _5192_/B _5087_/B _5250_/D _5127_/A vssd1 vssd1 vccd1 vccd1 _5202_/A sky130_fd_sc_hd__or4_1
X_8915_ _8915_/A _4398_/Y vssd1 vssd1 vccd1 vccd1 io_out[2] sky130_fd_sc_hd__ebufn_8
XFILLER_71_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5989_ _6077_/A _6077_/B vssd1 vssd1 vccd1 vccd1 _6000_/A sky130_fd_sc_hd__xnor2_2
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8777_ _8778_/CLK _8777_/D vssd1 vssd1 vccd1 vccd1 _8777_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7728_ _8780_/Q _8656_/Q vssd1 vssd1 vccd1 vccd1 _7752_/B sky130_fd_sc_hd__xnor2_2
XFILLER_12_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7659_ _7775_/A _8767_/Q vssd1 vssd1 vccd1 vccd1 _7661_/A sky130_fd_sc_hd__nand2_1
XFILLER_97_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_3_4_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_9_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5010_ _5187_/A _5119_/A vssd1 vssd1 vccd1 vccd1 _5172_/C sky130_fd_sc_hd__or2_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6961_ _7400_/A _6961_/B vssd1 vssd1 vccd1 vccd1 _6967_/A sky130_fd_sc_hd__nor2_1
X_8700_ _8732_/CLK _8700_/D vssd1 vssd1 vccd1 vccd1 _8700_/Q sky130_fd_sc_hd__dfxtp_1
X_5912_ _5971_/A _5971_/B vssd1 vssd1 vccd1 vccd1 _5940_/A sky130_fd_sc_hd__xor2_1
X_6892_ _6892_/A _6892_/B vssd1 vssd1 vccd1 vccd1 _6892_/Y sky130_fd_sc_hd__nor2_1
XFILLER_34_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5843_ _5843_/A _5888_/B _5843_/C vssd1 vssd1 vccd1 vccd1 _5887_/A sky130_fd_sc_hd__nand3_1
X_8631_ _8730_/CLK _8631_/D vssd1 vssd1 vccd1 vccd1 _8631_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8562_ _8562_/A _8562_/B _8562_/C vssd1 vssd1 vccd1 vccd1 _8563_/B sky130_fd_sc_hd__and3_1
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5774_ _5769_/Y _5652_/B _5775_/A _5527_/A vssd1 vssd1 vccd1 vccd1 _5872_/A sky130_fd_sc_hd__o211a_2
X_7513_ _7513_/A _7513_/B vssd1 vssd1 vccd1 vccd1 _7514_/B sky130_fd_sc_hd__xor2_2
X_8493_ _8424_/A _8424_/B _8492_/X vssd1 vssd1 vccd1 vccd1 _8501_/A sky130_fd_sc_hd__a21oi_1
X_4725_ _5231_/A vssd1 vssd1 vccd1 vccd1 _5271_/A sky130_fd_sc_hd__clkbuf_2
X_4656_ _8643_/Q _4656_/B vssd1 vssd1 vccd1 vccd1 _4661_/C sky130_fd_sc_hd__and2_1
X_7444_ _7375_/B _7444_/B vssd1 vssd1 vccd1 vccd1 _7444_/X sky130_fd_sc_hd__and2b_1
X_4587_ _8681_/Q _4595_/B vssd1 vssd1 vccd1 vccd1 _4588_/A sky130_fd_sc_hd__and2_1
X_7375_ _7444_/B _7375_/B vssd1 vssd1 vccd1 vccd1 _7430_/A sky130_fd_sc_hd__xnor2_2
X_6326_ _6326_/A _6326_/B vssd1 vssd1 vccd1 vccd1 _6326_/Y sky130_fd_sc_hd__nor2_1
XFILLER_1_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6257_ _6257_/A _6257_/B vssd1 vssd1 vccd1 vccd1 _6284_/A sky130_fd_sc_hd__xnor2_1
XFILLER_88_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6188_ _6188_/A _6247_/A vssd1 vssd1 vccd1 vccd1 _6189_/B sky130_fd_sc_hd__xnor2_1
X_5208_ _5030_/Y _5207_/Y _5255_/A vssd1 vssd1 vccd1 vccd1 _5211_/C sky130_fd_sc_hd__a21oi_1
XFILLER_69_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5139_ _5139_/A vssd1 vssd1 vccd1 vccd1 _5197_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_29_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5490_ _6460_/A vssd1 vssd1 vccd1 vccd1 _7656_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_4510_ _8664_/Q vssd1 vssd1 vccd1 vccd1 _4878_/B sky130_fd_sc_hd__clkbuf_1
X_4441_ _4444_/A vssd1 vssd1 vccd1 vccd1 _4441_/Y sky130_fd_sc_hd__inv_2
X_7160_ _7332_/A vssd1 vssd1 vccd1 vccd1 _7434_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_98_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6111_ _5944_/Y _6251_/A _6016_/B _6019_/A _6019_/B vssd1 vssd1 vccd1 vccd1 _6156_/B
+ sky130_fd_sc_hd__a32o_1
X_4372_ _4376_/A vssd1 vssd1 vccd1 vccd1 _4372_/Y sky130_fd_sc_hd__inv_2
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7091_ _7092_/A _7092_/B _7093_/B vssd1 vssd1 vccd1 vccd1 _7096_/B sky130_fd_sc_hd__a21o_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6042_ _6042_/A _6042_/B vssd1 vssd1 vccd1 vccd1 _6043_/B sky130_fd_sc_hd__or2_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7993_ _7991_/B _8063_/A _8270_/B vssd1 vssd1 vccd1 vccd1 _7994_/C sky130_fd_sc_hd__a21o_1
XFILLER_81_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6944_ _7228_/A _7228_/B vssd1 vssd1 vccd1 vccd1 _7212_/A sky130_fd_sc_hd__xnor2_2
XFILLER_22_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8614_ _8606_/B _8614_/B vssd1 vssd1 vccd1 vccd1 _8615_/C sky130_fd_sc_hd__and2b_1
XFILLER_22_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6875_ _6875_/A _6875_/B vssd1 vssd1 vccd1 vccd1 _6922_/A sky130_fd_sc_hd__xnor2_2
X_5826_ _5826_/A vssd1 vssd1 vccd1 vccd1 _5980_/A sky130_fd_sc_hd__buf_2
XFILLER_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8545_ _8545_/A _8545_/B vssd1 vssd1 vccd1 vccd1 _8547_/C sky130_fd_sc_hd__xnor2_2
X_5757_ _5756_/A _5756_/B _5756_/C vssd1 vssd1 vccd1 vccd1 _5811_/C sky130_fd_sc_hd__a21o_1
XFILLER_22_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8476_ _8477_/A _8477_/B _8477_/C vssd1 vssd1 vccd1 vccd1 _8491_/A sky130_fd_sc_hd__o21ai_1
X_4708_ _5264_/A vssd1 vssd1 vccd1 vccd1 _5221_/A sky130_fd_sc_hd__clkbuf_2
X_5688_ _5688_/A vssd1 vssd1 vccd1 vccd1 _5991_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7427_ _7427_/A _7427_/B vssd1 vssd1 vccd1 vccd1 _7427_/Y sky130_fd_sc_hd__nand2_1
X_4639_ _4643_/C _4639_/B vssd1 vssd1 vccd1 vccd1 _8637_/D sky130_fd_sc_hd__nor2_1
X_7358_ _7320_/A _7320_/B _7319_/A vssd1 vssd1 vccd1 vccd1 _7374_/A sky130_fd_sc_hd__a21o_1
X_6309_ _6231_/A _6309_/B vssd1 vssd1 vccd1 vccd1 _6309_/X sky130_fd_sc_hd__and2b_1
X_7289_ _7192_/A _7192_/B _7288_/Y vssd1 vssd1 vccd1 vccd1 _7291_/B sky130_fd_sc_hd__a21oi_1
XFILLER_76_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4990_ _5269_/A _4995_/C _4989_/X vssd1 vssd1 vccd1 vccd1 _4990_/X sky130_fd_sc_hd__or3b_1
X_6660_ _6660_/A _6660_/B vssd1 vssd1 vccd1 vccd1 _6703_/B sky130_fd_sc_hd__and2_1
X_5611_ _5626_/A _5611_/B vssd1 vssd1 vccd1 vccd1 _5720_/B sky130_fd_sc_hd__xnor2_1
XFILLER_31_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6591_ _6590_/A _6597_/A _6590_/C vssd1 vssd1 vccd1 vccd1 _6591_/X sky130_fd_sc_hd__a21o_1
X_8330_ _8330_/A _8330_/B vssd1 vssd1 vccd1 vccd1 _8417_/A sky130_fd_sc_hd__or2_1
X_5542_ _5542_/A _5541_/Y vssd1 vssd1 vccd1 vccd1 _5554_/A sky130_fd_sc_hd__or2b_2
X_8261_ _8261_/A _8273_/B vssd1 vssd1 vccd1 vccd1 _8263_/B sky130_fd_sc_hd__nor2_1
X_5473_ _5472_/X _5467_/B _5465_/B vssd1 vssd1 vccd1 vccd1 _5475_/C sky130_fd_sc_hd__a21oi_1
X_8192_ _8122_/Y _8102_/B _8355_/A vssd1 vssd1 vccd1 vccd1 _8192_/Y sky130_fd_sc_hd__a21boi_1
X_7212_ _7212_/A _7230_/A vssd1 vssd1 vccd1 vccd1 _7213_/B sky130_fd_sc_hd__nand2_1
X_4424_ _4425_/A vssd1 vssd1 vccd1 vccd1 _4424_/Y sky130_fd_sc_hd__inv_2
X_7143_ _7147_/A _7147_/B _7142_/X vssd1 vssd1 vccd1 vccd1 _7146_/B sky130_fd_sc_hd__a21oi_1
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7074_ _7099_/A _7099_/B vssd1 vssd1 vccd1 vccd1 _7100_/A sky130_fd_sc_hd__nor2_1
XFILLER_86_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6025_ _6119_/A _6025_/B vssd1 vssd1 vccd1 vccd1 _6027_/B sky130_fd_sc_hd__nor2_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7976_ _7976_/A _7976_/B _7976_/C vssd1 vssd1 vccd1 vccd1 _7977_/B sky130_fd_sc_hd__and3_1
X_6927_ _7301_/A _7389_/A vssd1 vssd1 vccd1 vccd1 _6933_/A sky130_fd_sc_hd__nand2_1
X_6858_ _7378_/A _6858_/B _6858_/C vssd1 vssd1 vccd1 vccd1 _6861_/A sky130_fd_sc_hd__and3_1
X_5809_ _5804_/B _5809_/B vssd1 vssd1 vccd1 vccd1 _5881_/A sky130_fd_sc_hd__and2b_1
XFILLER_50_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8528_ _8528_/A _8528_/B vssd1 vssd1 vccd1 vccd1 _8528_/Y sky130_fd_sc_hd__nand2_1
XFILLER_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6789_ _7118_/A _6965_/A _7400_/B _6829_/A vssd1 vssd1 vccd1 vccd1 _6807_/A sky130_fd_sc_hd__and4_1
X_8459_ _8459_/A _8459_/B vssd1 vssd1 vccd1 vccd1 _8513_/A sky130_fd_sc_hd__nand2_1
XFILLER_89_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7830_ _8568_/C _7934_/B _8378_/B vssd1 vssd1 vccd1 vccd1 _7831_/B sky130_fd_sc_hd__nor3_1
X_7761_ _7761_/A _8568_/B vssd1 vssd1 vccd1 vccd1 _7773_/A sky130_fd_sc_hd__nand2_1
XFILLER_51_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4973_ _4973_/A _4973_/B vssd1 vssd1 vccd1 vccd1 _5224_/A sky130_fd_sc_hd__or2_1
XFILLER_17_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7692_ _8568_/A _7783_/A vssd1 vssd1 vccd1 vccd1 _7761_/A sky130_fd_sc_hd__nor2_1
X_6712_ _6694_/A _7050_/A _7392_/B _6707_/A vssd1 vssd1 vccd1 vccd1 _6713_/B sky130_fd_sc_hd__o22ai_1
XFILLER_32_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6643_ _7309_/A _7391_/A _6641_/X vssd1 vssd1 vccd1 vccd1 _6644_/B sky130_fd_sc_hd__a21o_1
X_6574_ _6570_/A _6567_/X _6569_/X _6573_/X vssd1 vssd1 vccd1 vccd1 _8749_/D sky130_fd_sc_hd__a22o_1
X_5525_ _5916_/A vssd1 vssd1 vccd1 vccd1 _5922_/A sky130_fd_sc_hd__clkbuf_2
X_8313_ _8315_/A _8315_/B vssd1 vssd1 vccd1 vccd1 _8562_/A sky130_fd_sc_hd__xnor2_1
X_8244_ _8244_/A _8244_/B vssd1 vssd1 vccd1 vccd1 _8245_/B sky130_fd_sc_hd__xnor2_1
X_5456_ _8706_/Q _5456_/B vssd1 vssd1 vccd1 vccd1 _5458_/A sky130_fd_sc_hd__and2b_1
X_4407_ _4407_/A vssd1 vssd1 vccd1 vccd1 _4407_/Y sky130_fd_sc_hd__inv_2
X_8175_ _8175_/A _8248_/C vssd1 vssd1 vccd1 vccd1 _8177_/B sky130_fd_sc_hd__xnor2_1
X_5387_ _8696_/Q _6528_/C _5387_/C vssd1 vssd1 vccd1 vccd1 _5395_/C sky130_fd_sc_hd__and3_1
XFILLER_99_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7126_ _7126_/A _7126_/B vssd1 vssd1 vccd1 vccd1 _7127_/B sky130_fd_sc_hd__nand2_1
XFILLER_101_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7057_ _7221_/A _7221_/B vssd1 vssd1 vccd1 vccd1 _7058_/B sky130_fd_sc_hd__xnor2_1
X_6008_ _6064_/A _6008_/B vssd1 vssd1 vccd1 vccd1 _6009_/B sky130_fd_sc_hd__nor2_1
XFILLER_74_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7959_ _7959_/A _7959_/B vssd1 vssd1 vccd1 vccd1 _7959_/Y sky130_fd_sc_hd__nor2_1
XFILLER_54_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8859__76 vssd1 vssd1 vccd1 vccd1 _8859__76/HI _8968_/A sky130_fd_sc_hd__conb_1
X_6290_ _6290_/A _6290_/B _6290_/C vssd1 vssd1 vccd1 vccd1 _6291_/B sky130_fd_sc_hd__or3_1
X_5310_ _8673_/Q _5313_/B vssd1 vssd1 vccd1 vccd1 _5310_/X sky130_fd_sc_hd__or2_1
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5241_ _5234_/X _5236_/X _5240_/X _4697_/B _4736_/A vssd1 vssd1 vccd1 vccd1 _5241_/X
+ sky130_fd_sc_hd__a221o_1
X_5172_ _5172_/A _5283_/B _5172_/C vssd1 vssd1 vccd1 vccd1 _5173_/B sky130_fd_sc_hd__or3_1
Xinput2 io_in[10] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__buf_2
X_8931_ _8931_/A _4418_/Y vssd1 vssd1 vccd1 vccd1 io_out[18] sky130_fd_sc_hd__ebufn_8
XFILLER_96_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7813_ _7813_/A _7813_/B _7813_/C vssd1 vssd1 vccd1 vccd1 _8155_/B sky130_fd_sc_hd__nand3_1
X_7744_ _7924_/A vssd1 vssd1 vccd1 vccd1 _8568_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4956_ _4956_/A vssd1 vssd1 vccd1 vccd1 _5224_/B sky130_fd_sc_hd__buf_2
X_7675_ _8769_/Q _8666_/Q vssd1 vssd1 vccd1 vccd1 _7708_/B sky130_fd_sc_hd__xnor2_4
XFILLER_32_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4887_ _4934_/A _4922_/A _5162_/A vssd1 vssd1 vccd1 vccd1 _4887_/X sky130_fd_sc_hd__o21a_1
X_6626_ _6768_/A vssd1 vssd1 vccd1 vccd1 _6898_/A sky130_fd_sc_hd__clkbuf_2
X_6557_ _6570_/A _8748_/Q _6588_/B _6628_/B _6583_/A vssd1 vssd1 vccd1 vccd1 _6557_/X
+ sky130_fd_sc_hd__a2111o_1
X_5508_ _7685_/A _8710_/Q vssd1 vssd1 vccd1 vccd1 _5508_/X sky130_fd_sc_hd__or2b_1
X_6488_ _6492_/C _6488_/B vssd1 vssd1 vccd1 vccd1 _8732_/D sky130_fd_sc_hd__nor2_1
X_8227_ _8227_/A vssd1 vssd1 vccd1 vccd1 _8552_/A sky130_fd_sc_hd__clkbuf_1
X_5439_ _5456_/B _5452_/A _5463_/B vssd1 vssd1 vccd1 vccd1 _5440_/D sky130_fd_sc_hd__o21a_1
X_8873__90 vssd1 vssd1 vccd1 vccd1 _8873__90/HI _8982_/A sky130_fd_sc_hd__conb_1
X_8158_ _8158_/A _8158_/B _8158_/C vssd1 vssd1 vccd1 vccd1 _8272_/A sky130_fd_sc_hd__and3_1
XFILLER_59_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7109_ _7117_/B _7117_/A vssd1 vssd1 vccd1 vccd1 _7111_/A sky130_fd_sc_hd__and2b_1
X_8089_ _7845_/A _7845_/B _7689_/A _7689_/B _7943_/Y vssd1 vssd1 vccd1 vccd1 _8330_/B
+ sky130_fd_sc_hd__a2111o_1
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_6_0_wb_clk_i clkbuf_4_7_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _8765_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4810_ _7589_/A _4810_/B _4810_/C vssd1 vssd1 vccd1 vccd1 _4811_/A sky130_fd_sc_hd__and3_1
XFILLER_92_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5790_ _5790_/A _5790_/B vssd1 vssd1 vccd1 vccd1 _5791_/B sky130_fd_sc_hd__and2_1
XFILLER_33_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4741_ _4741_/A _5301_/B vssd1 vssd1 vccd1 vccd1 _5296_/A sky130_fd_sc_hd__or2_1
X_4672_ _4674_/B _4672_/B _4672_/C vssd1 vssd1 vccd1 vccd1 _4673_/A sky130_fd_sc_hd__and3b_1
X_7460_ _7489_/A _6801_/C _7460_/S vssd1 vssd1 vccd1 vccd1 _7471_/A sky130_fd_sc_hd__mux2_1
X_6411_ _6413_/A _6413_/B vssd1 vssd1 vccd1 vccd1 _6411_/X sky130_fd_sc_hd__xor2_1
X_7391_ _7391_/A _7391_/B vssd1 vssd1 vccd1 vccd1 _7391_/Y sky130_fd_sc_hd__nor2_1
X_6342_ _6342_/A vssd1 vssd1 vccd1 vccd1 _6342_/Y sky130_fd_sc_hd__inv_2
X_6273_ _6193_/A _6275_/S _6194_/B _6274_/B vssd1 vssd1 vccd1 vccd1 _6276_/A sky130_fd_sc_hd__a22o_1
X_8012_ _8082_/A _8082_/B vssd1 vssd1 vccd1 vccd1 _8013_/B sky130_fd_sc_hd__xor2_1
X_5224_ _5224_/A _5224_/B _5224_/C _5224_/D vssd1 vssd1 vccd1 vccd1 _5224_/X sky130_fd_sc_hd__or4_1
XFILLER_96_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5155_ _5272_/B _5183_/A _5155_/C _5274_/B vssd1 vssd1 vccd1 vccd1 _5157_/D sky130_fd_sc_hd__or4_1
XFILLER_56_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5086_ _5086_/A vssd1 vssd1 vccd1 vccd1 _5127_/A sky130_fd_sc_hd__clkbuf_2
X_8914_ _8914_/A _4397_/Y vssd1 vssd1 vccd1 vccd1 io_out[1] sky130_fd_sc_hd__ebufn_8
XFILLER_25_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5988_ _5988_/A _5988_/B vssd1 vssd1 vccd1 vccd1 _6077_/B sky130_fd_sc_hd__xnor2_1
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8776_ _8776_/CLK _8776_/D vssd1 vssd1 vccd1 vccd1 _8776_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7727_ _7727_/A vssd1 vssd1 vccd1 vccd1 _7821_/A sky130_fd_sc_hd__clkbuf_2
X_4939_ _5108_/A _5041_/A vssd1 vssd1 vccd1 vccd1 _5201_/B sky130_fd_sc_hd__or2_2
X_7658_ _7665_/A _7651_/B _7666_/S vssd1 vssd1 vccd1 vccd1 _7662_/A sky130_fd_sc_hd__a21o_1
X_6609_ _8759_/Q vssd1 vssd1 vccd1 vccd1 _7558_/A sky130_fd_sc_hd__inv_2
XFILLER_20_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7589_ _7589_/A _7589_/B _7589_/C vssd1 vssd1 vccd1 vccd1 _7590_/A sky130_fd_sc_hd__and3_1
XFILLER_87_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8829__46 vssd1 vssd1 vccd1 vccd1 _8829__46/HI _8938_/A sky130_fd_sc_hd__conb_1
XFILLER_7_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6960_ _7123_/A _6960_/B vssd1 vssd1 vccd1 vccd1 _6961_/B sky130_fd_sc_hd__nand2_1
XFILLER_38_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5911_ _5911_/A _5911_/B vssd1 vssd1 vccd1 vccd1 _5971_/B sky130_fd_sc_hd__xor2_2
XFILLER_19_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6891_ _6891_/A _6891_/B vssd1 vssd1 vccd1 vccd1 _6982_/B sky130_fd_sc_hd__xor2_1
XFILLER_46_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5842_ _5888_/A _5841_/B _5841_/C vssd1 vssd1 vccd1 vccd1 _5843_/C sky130_fd_sc_hd__a21o_1
X_8630_ _7602_/A _8628_/Y _8629_/Y vssd1 vssd1 vccd1 vccd1 _8785_/D sky130_fd_sc_hd__a21oi_1
XFILLER_34_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5773_ _5773_/A _6165_/B vssd1 vssd1 vccd1 vccd1 _5775_/A sky130_fd_sc_hd__nor2_1
XFILLER_61_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8561_ _8561_/A _8561_/B vssd1 vssd1 vccd1 vccd1 _8561_/Y sky130_fd_sc_hd__nor2_1
XFILLER_21_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4724_ _4730_/A _4723_/X _4760_/A vssd1 vssd1 vccd1 vccd1 _8654_/D sky130_fd_sc_hd__a21boi_1
X_7512_ _7512_/A _7512_/B vssd1 vssd1 vccd1 vccd1 _7513_/B sky130_fd_sc_hd__xnor2_4
X_8492_ _8423_/A _8492_/B vssd1 vssd1 vccd1 vccd1 _8492_/X sky130_fd_sc_hd__and2b_1
X_4655_ _4655_/A vssd1 vssd1 vccd1 vccd1 _8642_/D sky130_fd_sc_hd__clkbuf_1
X_7443_ _7432_/A _7432_/B _7442_/Y vssd1 vssd1 vccd1 vccd1 _7512_/A sky130_fd_sc_hd__a21o_1
X_4586_ _5305_/A vssd1 vssd1 vccd1 vccd1 _4595_/B sky130_fd_sc_hd__clkbuf_2
X_7374_ _7374_/A _7374_/B vssd1 vssd1 vccd1 vccd1 _7375_/B sky130_fd_sc_hd__xnor2_1
XFILLER_89_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6325_ _6325_/A _6325_/B vssd1 vssd1 vccd1 vccd1 _6339_/A sky130_fd_sc_hd__xor2_1
X_6256_ _6256_/A _6256_/B vssd1 vssd1 vccd1 vccd1 _6257_/B sky130_fd_sc_hd__nor2_1
X_6187_ _6274_/A _6187_/B vssd1 vssd1 vccd1 vccd1 _6247_/A sky130_fd_sc_hd__xnor2_1
X_8843__60 vssd1 vssd1 vccd1 vccd1 _8843__60/HI _8952_/A sky130_fd_sc_hd__conb_1
X_5207_ _5209_/A _5207_/B vssd1 vssd1 vccd1 vccd1 _5207_/Y sky130_fd_sc_hd__nor2_1
X_5138_ _5138_/A _5280_/A vssd1 vssd1 vccd1 vccd1 _5139_/A sky130_fd_sc_hd__nand2_1
XFILLER_72_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5069_ _5281_/B _5228_/A _5069_/C _5069_/D vssd1 vssd1 vccd1 vccd1 _5069_/X sky130_fd_sc_hd__or4_1
XFILLER_25_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8759_ _8763_/CLK _8759_/D vssd1 vssd1 vccd1 vccd1 _8759_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4440_ _4444_/A vssd1 vssd1 vccd1 vccd1 _4440_/Y sky130_fd_sc_hd__inv_2
X_6110_ _6320_/A _6110_/B vssd1 vssd1 vccd1 vccd1 _6156_/A sky130_fd_sc_hd__xnor2_1
X_4371_ _4395_/A vssd1 vssd1 vccd1 vccd1 _4376_/A sky130_fd_sc_hd__clkbuf_2
X_7090_ _7090_/A _7090_/B vssd1 vssd1 vccd1 vccd1 _7093_/B sky130_fd_sc_hd__xnor2_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6041_ _6042_/A _6042_/B vssd1 vssd1 vccd1 vccd1 _6043_/A sky130_fd_sc_hd__nand2_1
XFILLER_100_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7992_ _8068_/A vssd1 vssd1 vccd1 vccd1 _8270_/B sky130_fd_sc_hd__clkbuf_2
X_6943_ _6943_/A vssd1 vssd1 vccd1 vccd1 _7228_/A sky130_fd_sc_hd__clkbuf_4
X_6874_ _7019_/A _6874_/B vssd1 vssd1 vccd1 vccd1 _6875_/B sky130_fd_sc_hd__xnor2_2
X_5825_ _6378_/C _5983_/A vssd1 vssd1 vccd1 vccd1 _5826_/A sky130_fd_sc_hd__or2_1
X_8613_ _8619_/A _8613_/B vssd1 vssd1 vccd1 vccd1 _8615_/B sky130_fd_sc_hd__or2_1
X_8544_ _8544_/A _8544_/B vssd1 vssd1 vccd1 vccd1 _8545_/B sky130_fd_sc_hd__xnor2_2
X_5756_ _5756_/A _5756_/B _5756_/C vssd1 vssd1 vccd1 vccd1 _5811_/B sky130_fd_sc_hd__nand3_1
X_8475_ _8475_/A _8475_/B vssd1 vssd1 vccd1 vccd1 _8477_/C sky130_fd_sc_hd__xor2_1
X_5687_ _5687_/A vssd1 vssd1 vccd1 vccd1 _6071_/A sky130_fd_sc_hd__buf_2
X_4707_ _8653_/Q vssd1 vssd1 vccd1 vccd1 _5264_/A sky130_fd_sc_hd__inv_2
X_7426_ _7473_/A _7473_/B vssd1 vssd1 vccd1 vccd1 _7505_/A sky130_fd_sc_hd__xor2_2
X_4638_ _8637_/Q _4636_/A _4628_/X vssd1 vssd1 vccd1 vccd1 _4639_/B sky130_fd_sc_hd__o21ai_1
X_7357_ _7484_/S _7339_/B _7356_/X vssd1 vssd1 vccd1 vccd1 _7444_/B sky130_fd_sc_hd__a21o_1
X_4569_ _8671_/Q vssd1 vssd1 vccd1 vccd1 _4814_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6308_ _6234_/A _6234_/B _6307_/X vssd1 vssd1 vccd1 vccd1 _6315_/A sky130_fd_sc_hd__a21oi_1
X_7288_ _7288_/A _7288_/B vssd1 vssd1 vccd1 vccd1 _7288_/Y sky130_fd_sc_hd__nor2_1
X_6239_ _6343_/B _6239_/B vssd1 vssd1 vccd1 vccd1 _6242_/A sky130_fd_sc_hd__xnor2_1
XFILLER_103_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5610_ _5725_/A _5892_/A _5594_/A _5609_/Y vssd1 vssd1 vccd1 vccd1 _5611_/B sky130_fd_sc_hd__o211a_1
X_6590_ _6590_/A _6597_/A _6590_/C vssd1 vssd1 vccd1 vccd1 _6602_/A sky130_fd_sc_hd__nand3_1
X_5541_ _8712_/Q _7775_/B vssd1 vssd1 vccd1 vccd1 _5541_/Y sky130_fd_sc_hd__nand2_1
XFILLER_31_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8260_ _8248_/B _8158_/B _8158_/C vssd1 vssd1 vccd1 vccd1 _8266_/A sky130_fd_sc_hd__a21bo_1
X_5472_ _5478_/B _5463_/B vssd1 vssd1 vccd1 vccd1 _5472_/X sky130_fd_sc_hd__or2b_1
X_7211_ _7331_/A vssd1 vssd1 vccd1 vccd1 _7230_/A sky130_fd_sc_hd__inv_2
X_4423_ _4425_/A vssd1 vssd1 vccd1 vccd1 _4423_/Y sky130_fd_sc_hd__inv_2
X_8191_ _8355_/B vssd1 vssd1 vccd1 vccd1 _8418_/A sky130_fd_sc_hd__clkbuf_2
X_7142_ _7141_/A _7142_/B vssd1 vssd1 vccd1 vccd1 _7142_/X sky130_fd_sc_hd__and2b_1
XFILLER_98_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7073_ _7080_/D _7073_/B vssd1 vssd1 vccd1 vccd1 _7099_/B sky130_fd_sc_hd__xnor2_1
XFILLER_100_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6024_ _6024_/A _6024_/B vssd1 vssd1 vccd1 vccd1 _6025_/B sky130_fd_sc_hd__nor2_1
X_8813__30 vssd1 vssd1 vccd1 vccd1 _8813__30/HI _8908_/A sky130_fd_sc_hd__conb_1
XFILLER_58_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7975_ _7976_/A _7976_/B _7976_/C vssd1 vssd1 vccd1 vccd1 _8053_/A sky130_fd_sc_hd__a21oi_1
XFILLER_54_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6926_ _6799_/A _7389_/A _7231_/A vssd1 vssd1 vccd1 vccd1 _7228_/B sky130_fd_sc_hd__o21a_2
XFILLER_54_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6857_ _6999_/A _6857_/B vssd1 vssd1 vccd1 vccd1 _6858_/C sky130_fd_sc_hd__and2_1
X_5808_ _5709_/Y _6394_/A _5807_/X vssd1 vssd1 vccd1 vccd1 _6390_/A sky130_fd_sc_hd__a21oi_1
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6788_ _6788_/A _6788_/B vssd1 vssd1 vccd1 vccd1 _6829_/A sky130_fd_sc_hd__xnor2_2
X_8527_ _8527_/A _8527_/B vssd1 vssd1 vccd1 vccd1 _8533_/A sky130_fd_sc_hd__nor2_1
XFILLER_6_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5739_ _6433_/A _6673_/B vssd1 vssd1 vccd1 vccd1 _5739_/Y sky130_fd_sc_hd__nand2_1
X_8458_ _8394_/A _8394_/B _8394_/C _8457_/X vssd1 vssd1 vccd1 vccd1 _8521_/A sky130_fd_sc_hd__a31o_1
XFILLER_89_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8389_ _8389_/A _8389_/B vssd1 vssd1 vccd1 vccd1 _8463_/B sky130_fd_sc_hd__nor2_1
X_7409_ _7409_/A _7409_/B vssd1 vssd1 vccd1 vccd1 _7410_/B sky130_fd_sc_hd__nand2_1
XFILLER_89_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7760_ _7867_/A _7760_/B vssd1 vssd1 vccd1 vccd1 _7772_/A sky130_fd_sc_hd__nand2_1
X_4972_ _5170_/A _4972_/B _4972_/C vssd1 vssd1 vccd1 vccd1 _4972_/X sky130_fd_sc_hd__or3_1
X_7691_ _8024_/A _7854_/A vssd1 vssd1 vccd1 vccd1 _7783_/A sky130_fd_sc_hd__nand2_1
X_6711_ _6924_/A _6725_/A vssd1 vssd1 vccd1 vccd1 _6713_/A sky130_fd_sc_hd__or2_1
XFILLER_32_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6642_ _7120_/A _6641_/X vssd1 vssd1 vccd1 vccd1 _6644_/A sky130_fd_sc_hd__or2b_1
XFILLER_32_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8312_ _8312_/A _8312_/B vssd1 vssd1 vccd1 vccd1 _8315_/B sky130_fd_sc_hd__xnor2_1
X_6573_ _6571_/Y _6573_/B vssd1 vssd1 vccd1 vccd1 _6573_/X sky130_fd_sc_hd__and2b_1
X_5524_ _5531_/D vssd1 vssd1 vccd1 vccd1 _5861_/B sky130_fd_sc_hd__clkbuf_2
X_8243_ _8363_/A _8243_/B vssd1 vssd1 vccd1 vccd1 _8244_/B sky130_fd_sc_hd__nor2_1
X_5455_ _5452_/A _5449_/X _5450_/X _5454_/Y vssd1 vssd1 vccd1 vccd1 _8708_/D sky130_fd_sc_hd__a22o_1
X_4406_ _4407_/A vssd1 vssd1 vccd1 vccd1 _4406_/Y sky130_fd_sc_hd__clkinv_4
X_8174_ _8258_/A _8258_/B vssd1 vssd1 vccd1 vccd1 _8248_/C sky130_fd_sc_hd__xor2_1
X_7125_ _7125_/A vssd1 vssd1 vccd1 vccd1 _7128_/A sky130_fd_sc_hd__inv_2
X_5386_ _6528_/C _5387_/C _5385_/Y vssd1 vssd1 vccd1 vccd1 _8695_/D sky130_fd_sc_hd__a21oi_1
XFILLER_86_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7056_ _7056_/A _7056_/B vssd1 vssd1 vccd1 vccd1 _7221_/B sky130_fd_sc_hd__xor2_1
X_6007_ _6007_/A _6007_/B _6323_/A vssd1 vssd1 vccd1 vccd1 _6008_/B sky130_fd_sc_hd__and3_1
XFILLER_74_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7958_ _7958_/A _7958_/B vssd1 vssd1 vccd1 vccd1 _7962_/A sky130_fd_sc_hd__xnor2_1
XFILLER_15_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7889_ _7889_/A _7889_/B vssd1 vssd1 vccd1 vccd1 _7890_/A sky130_fd_sc_hd__and2_1
X_6909_ _6869_/B _6907_/Y _6909_/S vssd1 vssd1 vccd1 vccd1 _6914_/A sky130_fd_sc_hd__mux2_1
XFILLER_42_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5240_ _5237_/X _5238_/X _5239_/X vssd1 vssd1 vccd1 vccd1 _5240_/X sky130_fd_sc_hd__o21ba_1
XFILLER_68_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5171_ _5179_/B _5171_/B _5265_/B _5238_/B vssd1 vssd1 vccd1 vccd1 _5171_/X sky130_fd_sc_hd__or4_1
XFILLER_68_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8930_ _8930_/A _4417_/Y vssd1 vssd1 vccd1 vccd1 io_out[17] sky130_fd_sc_hd__ebufn_8
XFILLER_68_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7812_ _7913_/A _8381_/B _8155_/C vssd1 vssd1 vccd1 vccd1 _8010_/A sky130_fd_sc_hd__or3b_2
XFILLER_24_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7743_ _7902_/A vssd1 vssd1 vccd1 vccd1 _7924_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_24_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4955_ _4563_/X _4856_/Y _4946_/X _5136_/A _4954_/X vssd1 vssd1 vccd1 vccd1 _4955_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_51_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7674_ _7946_/A vssd1 vssd1 vccd1 vccd1 _8568_/A sky130_fd_sc_hd__clkbuf_2
X_4886_ _4934_/A _4921_/A _4889_/B _5032_/B _4885_/Y vssd1 vssd1 vccd1 vccd1 _5162_/A
+ sky130_fd_sc_hd__o221a_1
X_6625_ _6645_/A _6647_/B vssd1 vssd1 vccd1 vccd1 _6768_/A sky130_fd_sc_hd__xnor2_1
X_6556_ _8753_/Q vssd1 vssd1 vccd1 vccd1 _6758_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5507_ _8668_/Q vssd1 vssd1 vccd1 vccd1 _7685_/A sky130_fd_sc_hd__buf_2
X_8226_ _8312_/A _8312_/B vssd1 vssd1 vccd1 vccd1 _8227_/A sky130_fd_sc_hd__and2_1
X_6487_ _8732_/Q _6485_/A _6465_/X vssd1 vssd1 vccd1 vccd1 _6488_/B sky130_fd_sc_hd__o21ai_1
X_5438_ _5478_/B vssd1 vssd1 vccd1 vccd1 _5477_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_8157_ _8157_/A _8173_/B vssd1 vssd1 vccd1 vccd1 _8158_/C sky130_fd_sc_hd__nand2_1
XFILLER_87_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5369_ _8690_/Q _5372_/C vssd1 vssd1 vccd1 vccd1 _5371_/A sky130_fd_sc_hd__and2_1
XFILLER_101_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8088_ _8349_/A _8088_/B vssd1 vssd1 vccd1 vccd1 _8327_/A sky130_fd_sc_hd__nand2b_4
X_7108_ _7108_/A _7127_/A vssd1 vssd1 vccd1 vccd1 _7117_/A sky130_fd_sc_hd__nand2_1
XFILLER_87_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7039_ _7039_/A _7196_/A vssd1 vssd1 vccd1 vccd1 _7040_/B sky130_fd_sc_hd__xor2_1
XFILLER_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4740_ _4740_/A _4973_/A vssd1 vssd1 vccd1 vccd1 _5301_/B sky130_fd_sc_hd__nor2_1
XFILLER_14_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4671_ _8646_/Q _8647_/Q _4665_/B _8648_/Q vssd1 vssd1 vccd1 vccd1 _4672_/C sky130_fd_sc_hd__a31o_1
X_6410_ _6402_/S _6407_/B _6406_/A vssd1 vssd1 vccd1 vccd1 _6413_/B sky130_fd_sc_hd__o21ai_1
X_7390_ _7390_/A _7390_/B vssd1 vssd1 vccd1 vccd1 _7451_/A sky130_fd_sc_hd__xnor2_2
X_6341_ _6341_/A _6341_/B vssd1 vssd1 vccd1 vccd1 _6349_/A sky130_fd_sc_hd__xnor2_1
X_6272_ _6205_/A _6205_/B _6204_/A vssd1 vssd1 vccd1 vccd1 _6281_/A sky130_fd_sc_hd__a21o_1
X_8011_ _8376_/A _8011_/B vssd1 vssd1 vccd1 vccd1 _8082_/B sky130_fd_sc_hd__xnor2_1
X_5223_ _4995_/A _5250_/B _5221_/B _5217_/X _5222_/X vssd1 vssd1 vccd1 vccd1 _5224_/D
+ sky130_fd_sc_hd__o41a_1
XFILLER_102_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5154_ _5154_/A _5154_/B vssd1 vssd1 vccd1 vccd1 _5154_/X sky130_fd_sc_hd__or2_1
XFILLER_96_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5085_ _5085_/A vssd1 vssd1 vccd1 vccd1 _5192_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_29_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8913_ _8913_/A _4487_/Y vssd1 vssd1 vccd1 vccd1 io_out[0] sky130_fd_sc_hd__ebufn_8
XFILLER_56_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5987_ _6088_/A _6185_/A _6089_/A vssd1 vssd1 vccd1 vccd1 _5988_/B sky130_fd_sc_hd__o21a_1
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8775_ _8776_/CLK _8775_/D vssd1 vssd1 vccd1 vccd1 _8775_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7726_ _8655_/Q _8779_/Q vssd1 vssd1 vccd1 vccd1 _7727_/A sky130_fd_sc_hd__or2b_1
X_4938_ _4938_/A _5149_/B vssd1 vssd1 vccd1 vccd1 _5041_/A sky130_fd_sc_hd__or2_1
X_7657_ _7665_/A _6483_/X _7656_/X _7627_/X vssd1 vssd1 vccd1 vccd1 _8772_/D sky130_fd_sc_hd__a22o_1
X_4869_ _5108_/A vssd1 vssd1 vccd1 vccd1 _5209_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6608_ _7739_/B _8759_/Q vssd1 vssd1 vccd1 vccd1 _6648_/A sky130_fd_sc_hd__nand2b_2
X_7588_ _7587_/B _7587_/C _7587_/A vssd1 vssd1 vccd1 vccd1 _7589_/C sky130_fd_sc_hd__o21ai_1
X_6539_ _8760_/Q vssd1 vssd1 vccd1 vccd1 _7556_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_97_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8209_ _8325_/B _8497_/A vssd1 vssd1 vccd1 vccd1 _8236_/A sky130_fd_sc_hd__nor2_1
XFILLER_75_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5910_ _5897_/A _5907_/Y _6024_/A vssd1 vssd1 vccd1 vccd1 _5911_/B sky130_fd_sc_hd__a21oi_2
XFILLER_19_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6890_ _6892_/A _6892_/B vssd1 vssd1 vccd1 vccd1 _6982_/A sky130_fd_sc_hd__xor2_1
XFILLER_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5841_ _5888_/A _5841_/B _5841_/C vssd1 vssd1 vccd1 vccd1 _5888_/B sky130_fd_sc_hd__nand3_1
XFILLER_61_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5772_ _5853_/B vssd1 vssd1 vccd1 vccd1 _6165_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_8560_ _8559_/B _8559_/C _8559_/A vssd1 vssd1 vccd1 vccd1 _8561_/B sky130_fd_sc_hd__a21oi_1
X_8491_ _8491_/A _8491_/B vssd1 vssd1 vccd1 vccd1 _8545_/A sky130_fd_sc_hd__xnor2_1
X_4723_ _5271_/B _4745_/A vssd1 vssd1 vccd1 vccd1 _4723_/X sky130_fd_sc_hd__or2_1
X_7511_ _7511_/A _7511_/B vssd1 vssd1 vccd1 vccd1 _7512_/B sky130_fd_sc_hd__xnor2_2
X_7442_ _7442_/A _7442_/B vssd1 vssd1 vccd1 vccd1 _7442_/Y sky130_fd_sc_hd__nor2_1
X_4654_ _4656_/B _4672_/B _4654_/C vssd1 vssd1 vccd1 vccd1 _4655_/A sky130_fd_sc_hd__and3b_1
X_7373_ _7373_/A _7373_/B vssd1 vssd1 vccd1 vccd1 _7374_/B sky130_fd_sc_hd__xnor2_1
X_4585_ _4585_/A vssd1 vssd1 vccd1 vccd1 _8934_/A sky130_fd_sc_hd__clkbuf_1
X_6324_ _6264_/A _6264_/B _6265_/A _6323_/X vssd1 vssd1 vccd1 vccd1 _6325_/B sky130_fd_sc_hd__o31ai_1
XFILLER_88_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6255_ _6255_/A _6255_/B _6255_/C vssd1 vssd1 vccd1 vccd1 _6256_/B sky130_fd_sc_hd__and3_1
XFILLER_103_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5206_ _5206_/A _5206_/B vssd1 vssd1 vccd1 vccd1 _5207_/B sky130_fd_sc_hd__or2_1
X_6186_ _6186_/A _6186_/B vssd1 vssd1 vccd1 vccd1 _6187_/B sky130_fd_sc_hd__nor2_1
XFILLER_69_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5137_ _4964_/X _5250_/C _5250_/D _5149_/C _5136_/X vssd1 vssd1 vccd1 vccd1 _5137_/X
+ sky130_fd_sc_hd__o41a_1
XFILLER_84_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5068_ _5182_/A _5285_/A vssd1 vssd1 vccd1 vccd1 _5069_/D sky130_fd_sc_hd__or2_1
XFILLER_84_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8758_ _8758_/CLK _8758_/D vssd1 vssd1 vccd1 vccd1 _8758_/Q sky130_fd_sc_hd__dfxtp_1
X_7709_ _8025_/A vssd1 vssd1 vccd1 vccd1 _8325_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8689_ _8704_/CLK _8689_/D vssd1 vssd1 vccd1 vccd1 _8689_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4370_ input1/X vssd1 vssd1 vccd1 vccd1 _4395_/A sky130_fd_sc_hd__clkbuf_2
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6040_ _6121_/B _6040_/B vssd1 vssd1 vccd1 vccd1 _6042_/B sky130_fd_sc_hd__xnor2_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7991_ _8068_/A _7991_/B _8063_/A vssd1 vssd1 vccd1 vccd1 _8063_/B sky130_fd_sc_hd__nand3_1
X_6942_ _6881_/A _6881_/B _6887_/B _6888_/B _6888_/A vssd1 vssd1 vccd1 vccd1 _6994_/A
+ sky130_fd_sc_hd__a32o_1
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6873_ _6873_/A _6873_/B vssd1 vssd1 vccd1 vccd1 _6874_/B sky130_fd_sc_hd__or2_1
X_5824_ _6081_/A _5824_/B vssd1 vssd1 vccd1 vccd1 _5829_/A sky130_fd_sc_hd__nand2_1
X_8612_ _8626_/A _8612_/B vssd1 vssd1 vccd1 vccd1 _8613_/B sky130_fd_sc_hd__and2b_1
XFILLER_22_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8543_ _8543_/A _8543_/B vssd1 vssd1 vccd1 vccd1 _8544_/B sky130_fd_sc_hd__xnor2_1
X_5755_ _5845_/A _5755_/B vssd1 vssd1 vccd1 vccd1 _5756_/C sky130_fd_sc_hd__nor2_1
X_8474_ _8539_/A _8539_/B vssd1 vssd1 vccd1 vccd1 _8475_/B sky130_fd_sc_hd__xnor2_1
X_5686_ _5697_/A _5686_/B vssd1 vssd1 vccd1 vccd1 _5704_/A sky130_fd_sc_hd__nand2_1
X_4706_ _5136_/A _4771_/A _4732_/B _4705_/X vssd1 vssd1 vccd1 vccd1 _8652_/D sky130_fd_sc_hd__o211a_1
X_7425_ _7425_/A _7425_/B vssd1 vssd1 vccd1 vccd1 _7473_/B sky130_fd_sc_hd__xnor2_1
X_4637_ _8636_/Q _8637_/Q _4637_/C vssd1 vssd1 vccd1 vccd1 _4643_/C sky130_fd_sc_hd__and3_1
XFILLER_89_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7356_ _7338_/B _7356_/B vssd1 vssd1 vccd1 vccd1 _7356_/X sky130_fd_sc_hd__and2b_1
X_4568_ _4823_/A _4568_/B _4568_/C _4935_/A vssd1 vssd1 vccd1 vccd1 _4574_/C sky130_fd_sc_hd__or4_1
XFILLER_103_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6307_ _6233_/A _6307_/B vssd1 vssd1 vccd1 vccd1 _6307_/X sky130_fd_sc_hd__and2b_1
X_7287_ _7420_/A _7287_/B vssd1 vssd1 vccd1 vccd1 _7291_/A sky130_fd_sc_hd__xor2_1
X_4499_ _5249_/B _4740_/A vssd1 vssd1 vccd1 vccd1 _4565_/B sky130_fd_sc_hd__or2_1
XFILLER_103_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6238_ _6238_/A _6238_/B vssd1 vssd1 vccd1 vccd1 _6239_/B sky130_fd_sc_hd__xnor2_1
X_6169_ _6169_/A _6169_/B vssd1 vssd1 vccd1 vccd1 _6172_/A sky130_fd_sc_hd__or2_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5540_ _8712_/Q _7775_/B vssd1 vssd1 vccd1 vccd1 _5542_/A sky130_fd_sc_hd__nor2_1
X_5471_ _8711_/Q _5477_/B vssd1 vssd1 vccd1 vccd1 _5475_/B sky130_fd_sc_hd__or2b_1
XFILLER_8_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7210_ _7370_/A _7370_/B vssd1 vssd1 vccd1 vccd1 _7334_/A sky130_fd_sc_hd__nand2_1
X_4422_ _4425_/A vssd1 vssd1 vccd1 vccd1 _4422_/Y sky130_fd_sc_hd__inv_2
X_8190_ _8190_/A _8190_/B vssd1 vssd1 vccd1 vccd1 _8355_/B sky130_fd_sc_hd__or2_2
XFILLER_98_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7141_ _7141_/A _7142_/B vssd1 vssd1 vccd1 vccd1 _7147_/B sky130_fd_sc_hd__xnor2_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7072_ _7176_/A _7080_/C _6635_/A vssd1 vssd1 vccd1 vccd1 _7073_/B sky130_fd_sc_hd__a21o_1
X_6023_ _6024_/A _6024_/B vssd1 vssd1 vccd1 vccd1 _6119_/A sky130_fd_sc_hd__and2_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7974_ _7974_/A _7974_/B vssd1 vssd1 vccd1 vccd1 _7976_/C sky130_fd_sc_hd__or2_1
X_6925_ _6925_/A vssd1 vssd1 vccd1 vccd1 _7231_/A sky130_fd_sc_hd__clkbuf_2
X_6856_ _6856_/A _7182_/A vssd1 vssd1 vccd1 vccd1 _6857_/B sky130_fd_sc_hd__nand2_1
X_5807_ _5962_/B _5807_/B vssd1 vssd1 vccd1 vccd1 _5807_/X sky130_fd_sc_hd__xor2_1
XFILLER_50_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6787_ _6801_/B _6787_/B vssd1 vssd1 vccd1 vccd1 _6788_/B sky130_fd_sc_hd__and2_1
X_8526_ _8526_/A _8526_/B vssd1 vssd1 vccd1 vccd1 _8534_/A sky130_fd_sc_hd__xnor2_1
X_5738_ _5749_/A _5993_/B vssd1 vssd1 vccd1 vccd1 _5827_/A sky130_fd_sc_hd__nor2_1
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8457_ _8393_/A _8457_/B vssd1 vssd1 vccd1 vccd1 _8457_/X sky130_fd_sc_hd__and2b_1
X_5669_ _5670_/A _5670_/B vssd1 vssd1 vccd1 vccd1 _5799_/A sky130_fd_sc_hd__or2_1
X_8388_ _8387_/A _8387_/B _8387_/C vssd1 vssd1 vccd1 vccd1 _8394_/B sky130_fd_sc_hd__a21o_1
X_7408_ _7457_/B _7408_/B vssd1 vssd1 vccd1 vccd1 _7410_/A sky130_fd_sc_hd__xnor2_1
X_7339_ _7373_/A _7339_/B vssd1 vssd1 vccd1 vccd1 _7340_/B sky130_fd_sc_hd__xnor2_2
XFILLER_1_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_2_1_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_68_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4971_ _4563_/X _4953_/X _4856_/Y _4950_/X _4555_/X vssd1 vssd1 vccd1 vccd1 _4972_/C
+ sky130_fd_sc_hd__o221a_1
X_7690_ _8092_/A vssd1 vssd1 vccd1 vccd1 _7854_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_17_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6710_ _7302_/B _7002_/C vssd1 vssd1 vccd1 vccd1 _6725_/A sky130_fd_sc_hd__or2_1
XFILLER_32_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6641_ _7141_/A _7186_/B _6641_/C vssd1 vssd1 vccd1 vccd1 _6641_/X sky130_fd_sc_hd__and3_1
X_8311_ _8311_/A _8311_/B vssd1 vssd1 vccd1 vccd1 _8315_/A sky130_fd_sc_hd__nand2_1
X_6572_ _6621_/A _6572_/B vssd1 vssd1 vccd1 vccd1 _6573_/B sky130_fd_sc_hd__nand2_1
X_5523_ _6169_/A vssd1 vssd1 vccd1 vccd1 _5531_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_8242_ _8527_/A _8242_/B vssd1 vssd1 vccd1 vccd1 _8243_/B sky130_fd_sc_hd__and2_1
X_5454_ _8707_/Q _5454_/B vssd1 vssd1 vccd1 vccd1 _5454_/Y sky130_fd_sc_hd__xnor2_1
X_4405_ _4407_/A vssd1 vssd1 vccd1 vccd1 _4405_/Y sky130_fd_sc_hd__inv_2
X_8173_ _8264_/A _8173_/B vssd1 vssd1 vccd1 vccd1 _8258_/B sky130_fd_sc_hd__xor2_1
X_5385_ _6528_/C _5387_/C _5409_/A vssd1 vssd1 vccd1 vccd1 _5385_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_99_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7124_ _7119_/X _7140_/B _7139_/A vssd1 vssd1 vccd1 vccd1 _7125_/A sky130_fd_sc_hd__a21o_1
X_7055_ _7120_/B _7181_/B vssd1 vssd1 vccd1 vccd1 _7056_/B sky130_fd_sc_hd__or2_1
XFILLER_101_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6006_ _6007_/A _6007_/B _6323_/A vssd1 vssd1 vccd1 vccd1 _6064_/A sky130_fd_sc_hd__a21oi_2
XFILLER_55_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7957_ _8023_/B _7957_/B vssd1 vssd1 vccd1 vccd1 _7958_/B sky130_fd_sc_hd__xnor2_1
X_7888_ _7888_/A _7888_/B vssd1 vssd1 vccd1 vccd1 _7889_/B sky130_fd_sc_hd__or2_1
X_6908_ _7262_/B _7080_/C vssd1 vssd1 vccd1 vccd1 _6909_/S sky130_fd_sc_hd__nor2_1
XFILLER_50_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6839_ _6840_/A _6840_/B vssd1 vssd1 vccd1 vccd1 _6839_/X sky130_fd_sc_hd__or2_1
X_8509_ _8509_/A _8509_/B vssd1 vssd1 vccd1 vccd1 _8510_/B sky130_fd_sc_hd__xor2_1
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5170_ _5170_/A _5170_/B _5170_/C vssd1 vssd1 vccd1 vccd1 _5170_/X sky130_fd_sc_hd__or3_1
XFILLER_96_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7811_ _7813_/A _7813_/C _7813_/B vssd1 vssd1 vccd1 vccd1 _8155_/C sky130_fd_sc_hd__a21o_1
XFILLER_64_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7742_ _7821_/A _7752_/B vssd1 vssd1 vccd1 vccd1 _7902_/A sky130_fd_sc_hd__xor2_1
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4954_ _4702_/D _5209_/B _4995_/C _4950_/X _4953_/X vssd1 vssd1 vccd1 vccd1 _4954_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_20_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7673_ _7762_/A _7762_/B vssd1 vssd1 vccd1 vccd1 _7946_/A sky130_fd_sc_hd__and2_2
X_4885_ _5261_/B _5291_/A vssd1 vssd1 vccd1 vccd1 _4885_/Y sky130_fd_sc_hd__nor2_1
X_6624_ _8749_/Q _6630_/B vssd1 vssd1 vccd1 vccd1 _6647_/B sky130_fd_sc_hd__xnor2_2
X_6555_ _6593_/A _6560_/A _6552_/X _6588_/B vssd1 vssd1 vccd1 vccd1 _6555_/X sky130_fd_sc_hd__o31a_1
X_5506_ _8710_/Q _7684_/B vssd1 vssd1 vccd1 vccd1 _5509_/A sky130_fd_sc_hd__and2b_1
X_8225_ _8228_/A _8225_/B vssd1 vssd1 vccd1 vccd1 _8312_/B sky130_fd_sc_hd__xnor2_1
X_6486_ _8731_/Q _8732_/Q _6486_/C vssd1 vssd1 vccd1 vccd1 _6492_/C sky130_fd_sc_hd__and3_1
X_5437_ _8706_/Q vssd1 vssd1 vccd1 vccd1 _5478_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_8156_ _8157_/A _8173_/B vssd1 vssd1 vccd1 vccd1 _8158_/B sky130_fd_sc_hd__or2_1
XFILLER_87_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5368_ _5368_/A vssd1 vssd1 vccd1 vccd1 _8689_/D sky130_fd_sc_hd__clkbuf_1
X_8087_ _8147_/A _8147_/B vssd1 vssd1 vccd1 vccd1 _8117_/A sky130_fd_sc_hd__xor2_1
XFILLER_59_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7107_ _7126_/A _7126_/B vssd1 vssd1 vccd1 vccd1 _7127_/A sky130_fd_sc_hd__or2_1
X_5299_ _4558_/X _4716_/A _4744_/A _4555_/X vssd1 vssd1 vccd1 vccd1 _5300_/C sky130_fd_sc_hd__o211a_1
XFILLER_59_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7038_ _7038_/A _7038_/B vssd1 vssd1 vccd1 vccd1 _7196_/A sky130_fd_sc_hd__xnor2_1
XFILLER_55_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8864__81 vssd1 vssd1 vccd1 vccd1 _8864__81/HI _8973_/A sky130_fd_sc_hd__conb_1
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4670_ _8648_/Q _8647_/Q _4670_/C vssd1 vssd1 vccd1 vccd1 _4674_/B sky130_fd_sc_hd__and3_1
XFILLER_14_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6340_ _6340_/A _6340_/B vssd1 vssd1 vccd1 vccd1 _6341_/B sky130_fd_sc_hd__xnor2_1
XFILLER_6_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6271_ _6271_/A _6271_/B vssd1 vssd1 vccd1 vccd1 _6326_/A sky130_fd_sc_hd__xnor2_2
X_8010_ _8010_/A _8068_/A vssd1 vssd1 vccd1 vccd1 _8011_/B sky130_fd_sc_hd__xnor2_1
X_5222_ _5219_/X _5221_/X _5259_/C _5163_/B vssd1 vssd1 vccd1 vccd1 _5222_/X sky130_fd_sc_hd__a211o_1
X_5153_ _5159_/B _5225_/B _5153_/C _5156_/B vssd1 vssd1 vccd1 vccd1 _5154_/B sky130_fd_sc_hd__or4_1
XFILLER_96_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5084_ _5288_/A _5228_/C _5188_/B _5182_/A _5156_/B vssd1 vssd1 vccd1 vccd1 _5084_/X
+ sky130_fd_sc_hd__a2111o_1
X_8912_ _8912_/A _4396_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[31] sky130_fd_sc_hd__ebufn_8
XFILLER_84_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5986_ _5986_/A _5986_/B vssd1 vssd1 vccd1 vccd1 _6089_/A sky130_fd_sc_hd__nand2_1
X_8774_ _8785_/CLK _8774_/D vssd1 vssd1 vccd1 vccd1 _8774_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7725_ _7725_/A _7725_/B vssd1 vssd1 vccd1 vccd1 _7788_/A sky130_fd_sc_hd__nor2_4
X_4937_ _5108_/B _4937_/B vssd1 vssd1 vccd1 vccd1 _5149_/B sky130_fd_sc_hd__or2_2
X_7656_ _7666_/S _7656_/B _7656_/C vssd1 vssd1 vccd1 vccd1 _7656_/X sky130_fd_sc_hd__and3b_1
X_4868_ _5123_/A _5048_/A vssd1 vssd1 vccd1 vccd1 _5108_/A sky130_fd_sc_hd__or2_1
XFILLER_20_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6607_ _6607_/A vssd1 vssd1 vccd1 vccd1 _8754_/D sky130_fd_sc_hd__clkbuf_1
X_4799_ _4804_/B _4804_/C vssd1 vssd1 vccd1 vccd1 _4801_/B sky130_fd_sc_hd__or2_1
X_7587_ _7587_/A _7587_/B _7587_/C vssd1 vssd1 vccd1 vccd1 _7589_/B sky130_fd_sc_hd__or3_1
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6538_ _8761_/Q vssd1 vssd1 vccd1 vccd1 _7562_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6469_ _8726_/Q _6455_/B _8727_/Q vssd1 vssd1 vccd1 vccd1 _6470_/B sky130_fd_sc_hd__a21o_1
X_8208_ _8115_/A _8115_/B _8116_/A vssd1 vssd1 vccd1 vccd1 _8220_/A sky130_fd_sc_hd__a21oi_1
X_8139_ _8139_/A _8139_/B vssd1 vssd1 vccd1 vccd1 _8559_/A sky130_fd_sc_hd__nor2_1
XFILLER_101_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5840_ _5908_/A _5840_/B vssd1 vssd1 vccd1 vccd1 _5841_/C sky130_fd_sc_hd__xnor2_1
XFILLER_61_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5771_ _5650_/B _5652_/B _5770_/Y vssd1 vssd1 vccd1 vccd1 _5853_/B sky130_fd_sc_hd__a21o_1
XFILLER_61_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8490_ _8490_/A _8490_/B vssd1 vssd1 vccd1 vccd1 _8491_/B sky130_fd_sc_hd__xnor2_1
X_4722_ _5271_/B _4745_/A vssd1 vssd1 vccd1 vccd1 _4730_/A sky130_fd_sc_hd__nand2_1
X_7510_ _7510_/A _7510_/B vssd1 vssd1 vccd1 vccd1 _7511_/B sky130_fd_sc_hd__xnor2_1
X_7441_ _7434_/A _7434_/B _7433_/B _7433_/A vssd1 vssd1 vccd1 vccd1 _7513_/A sky130_fd_sc_hd__a2bb2o_1
X_4653_ _8640_/Q _8641_/Q _4647_/B _8642_/Q vssd1 vssd1 vccd1 vccd1 _4654_/C sky130_fd_sc_hd__a31o_1
X_4584_ _8680_/Q _4584_/B vssd1 vssd1 vccd1 vccd1 _4585_/A sky130_fd_sc_hd__and2_1
X_7372_ _7482_/B _7483_/B vssd1 vssd1 vccd1 vccd1 _7373_/B sky130_fd_sc_hd__xnor2_1
X_6323_ _6323_/A _6266_/B vssd1 vssd1 vccd1 vccd1 _6323_/X sky130_fd_sc_hd__or2b_1
X_6254_ _6255_/A _6255_/B _6255_/C vssd1 vssd1 vccd1 vccd1 _6256_/A sky130_fd_sc_hd__a21oi_1
XFILLER_103_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5205_ _4969_/X _5038_/A _4563_/X vssd1 vssd1 vccd1 vccd1 _5205_/X sky130_fd_sc_hd__o21a_1
X_6185_ _6185_/A _6185_/B _6185_/C vssd1 vssd1 vccd1 vccd1 _6186_/B sky130_fd_sc_hd__nor3_1
XFILLER_57_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5136_ _5136_/A _5136_/B _5136_/C _5251_/C vssd1 vssd1 vccd1 vccd1 _5136_/X sky130_fd_sc_hd__or4_1
XFILLER_57_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5067_ _5066_/A _5155_/C _5211_/B _5066_/Y _5272_/B vssd1 vssd1 vccd1 vccd1 _5069_/C
+ sky130_fd_sc_hd__o32a_1
XFILLER_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5969_ _5941_/B _5969_/B vssd1 vssd1 vccd1 vccd1 _5969_/X sky130_fd_sc_hd__and2b_1
XFILLER_40_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8757_ _8758_/CLK _8757_/D vssd1 vssd1 vccd1 vccd1 _8757_/Q sky130_fd_sc_hd__dfxtp_1
X_7708_ _7762_/A _7708_/B vssd1 vssd1 vccd1 vccd1 _8025_/A sky130_fd_sc_hd__xnor2_2
XFILLER_8_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8688_ _8704_/CLK _8688_/D vssd1 vssd1 vccd1 vccd1 _8688_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7639_ _7630_/A _7637_/B _7631_/Y vssd1 vssd1 vccd1 vccd1 _7640_/B sky130_fd_sc_hd__a21oi_1
XFILLER_4_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8834__51 vssd1 vssd1 vccd1 vccd1 _8834__51/HI _8943_/A sky130_fd_sc_hd__conb_1
XFILLER_57_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7990_ _8165_/C _8514_/A _8381_/B _7828_/B vssd1 vssd1 vccd1 vccd1 _8063_/A sky130_fd_sc_hd__or4b_1
XFILLER_81_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6941_ _6941_/A _6996_/B vssd1 vssd1 vccd1 vccd1 _6954_/A sky130_fd_sc_hd__xnor2_1
X_6872_ _7011_/A vssd1 vssd1 vccd1 vccd1 _7019_/A sky130_fd_sc_hd__buf_4
XFILLER_34_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5823_ _5890_/B _5822_/C _5822_/A vssd1 vssd1 vccd1 vccd1 _5830_/B sky130_fd_sc_hd__a21o_1
X_8611_ _8612_/B _8626_/A vssd1 vssd1 vccd1 vccd1 _8619_/A sky130_fd_sc_hd__and2b_1
XFILLER_34_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8542_ _8542_/A _8542_/B vssd1 vssd1 vccd1 vccd1 _8543_/B sky130_fd_sc_hd__xnor2_1
XFILLER_34_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5754_ _5754_/A _5754_/B _5754_/C vssd1 vssd1 vccd1 vccd1 _5755_/B sky130_fd_sc_hd__nor3_1
X_8473_ _8473_/A _8488_/B vssd1 vssd1 vccd1 vccd1 _8539_/B sky130_fd_sc_hd__xnor2_1
X_5685_ _5766_/A _5533_/A _6149_/C _5684_/Y vssd1 vssd1 vccd1 vccd1 _5686_/B sky130_fd_sc_hd__a31o_1
X_4705_ _4760_/A vssd1 vssd1 vccd1 vccd1 _4705_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7424_ _7293_/A _7292_/B _7290_/Y vssd1 vssd1 vccd1 vccd1 _7425_/B sky130_fd_sc_hd__a21oi_1
X_4636_ _4636_/A _4636_/B vssd1 vssd1 vccd1 vccd1 _8636_/D sky130_fd_sc_hd__nor2_1
X_7355_ _7342_/A _7342_/B _7354_/X vssd1 vssd1 vccd1 vccd1 _7442_/A sky130_fd_sc_hd__a21oi_4
X_6306_ _6238_/A _6238_/B _6305_/X vssd1 vssd1 vccd1 vccd1 _6316_/A sky130_fd_sc_hd__a21o_1
X_4567_ _4877_/B _4762_/A _4872_/B _4877_/A vssd1 vssd1 vccd1 vccd1 _4935_/A sky130_fd_sc_hd__or4bb_2
X_4498_ _6615_/B vssd1 vssd1 vccd1 vccd1 _4740_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7286_ _7416_/B _7286_/B vssd1 vssd1 vccd1 vccd1 _7287_/B sky130_fd_sc_hd__xor2_1
X_6237_ _6237_/A _6305_/B vssd1 vssd1 vccd1 vccd1 _6238_/B sky130_fd_sc_hd__xnor2_1
X_6168_ _6228_/A _6168_/B vssd1 vssd1 vccd1 vccd1 _6175_/A sky130_fd_sc_hd__xnor2_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5119_ _5119_/A _5119_/B vssd1 vssd1 vccd1 vccd1 _5197_/C sky130_fd_sc_hd__or2_1
XFILLER_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6099_ _6099_/A _6099_/B vssd1 vssd1 vccd1 vccd1 _6100_/B sky130_fd_sc_hd__nand2_1
XFILLER_17_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_3_3_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_7_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_25_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5470_ _5477_/B _5484_/A vssd1 vssd1 vccd1 vccd1 _5480_/A sky130_fd_sc_hd__or2b_1
XFILLER_8_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4421_ _4425_/A vssd1 vssd1 vccd1 vccd1 _4421_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7140_ _7140_/A _7140_/B vssd1 vssd1 vccd1 vccd1 _7142_/B sky130_fd_sc_hd__xnor2_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7071_ _6965_/A _6961_/B _6967_/A vssd1 vssd1 vccd1 vccd1 _7099_/A sky130_fd_sc_hd__a21o_1
X_6022_ _6057_/A _6058_/A vssd1 vssd1 vccd1 vccd1 _6024_/B sky130_fd_sc_hd__xnor2_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7973_ _7972_/A _7972_/B _7972_/C vssd1 vssd1 vccd1 vccd1 _7974_/B sky130_fd_sc_hd__o21a_1
XFILLER_39_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6924_ _6924_/A _7391_/B vssd1 vssd1 vccd1 vccd1 _6925_/A sky130_fd_sc_hd__or2_1
XFILLER_35_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6855_ _6856_/A _7182_/A vssd1 vssd1 vccd1 vccd1 _6999_/A sky130_fd_sc_hd__or2_1
XFILLER_22_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5806_ _5959_/A _5962_/A vssd1 vssd1 vccd1 vccd1 _5807_/B sky130_fd_sc_hd__nand2_1
XFILLER_22_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6786_ _6786_/A _6786_/B vssd1 vssd1 vccd1 vccd1 _6787_/B sky130_fd_sc_hd__or2_1
X_8525_ _8525_/A _8525_/B vssd1 vssd1 vccd1 vccd1 _8526_/B sky130_fd_sc_hd__xnor2_2
X_5737_ _5983_/A vssd1 vssd1 vccd1 vccd1 _5993_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_10_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8456_ _8456_/A _8456_/B vssd1 vssd1 vccd1 vccd1 _8467_/A sky130_fd_sc_hd__xor2_2
XFILLER_13_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5668_ _5531_/X _5556_/Y _5787_/B vssd1 vssd1 vccd1 vccd1 _5670_/B sky130_fd_sc_hd__a21bo_1
X_7407_ _7282_/A _7282_/B _7406_/X vssd1 vssd1 vccd1 vccd1 _7408_/B sky130_fd_sc_hd__o21a_1
X_8387_ _8387_/A _8387_/B _8387_/C vssd1 vssd1 vccd1 vccd1 _8394_/A sky130_fd_sc_hd__nand3_1
X_5599_ _5979_/A vssd1 vssd1 vccd1 vccd1 _6068_/A sky130_fd_sc_hd__clkbuf_2
X_4619_ _8632_/Q _8631_/Q vssd1 vssd1 vccd1 vccd1 _4620_/C sky130_fd_sc_hd__nand2_1
X_7338_ _7356_/B _7338_/B vssd1 vssd1 vccd1 vccd1 _7339_/B sky130_fd_sc_hd__xnor2_1
XFILLER_104_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7269_ _7268_/B _7268_/C _7268_/A vssd1 vssd1 vccd1 vccd1 _7270_/C sky130_fd_sc_hd__a21o_1
XFILLER_89_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8804__21 vssd1 vssd1 vccd1 vccd1 _8804__21/HI _8899_/A sky130_fd_sc_hd__conb_1
XFILLER_73_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4970_ _4946_/X _4965_/X _4967_/X _4969_/X _4558_/X vssd1 vssd1 vccd1 vccd1 _4972_/B
+ sky130_fd_sc_hd__o221a_1
X_6640_ _6647_/B _6707_/A _6793_/A vssd1 vssd1 vccd1 vccd1 _6641_/C sky130_fd_sc_hd__o21ai_1
X_6571_ _6621_/A _6572_/B vssd1 vssd1 vccd1 vccd1 _6571_/Y sky130_fd_sc_hd__nor2_1
X_5522_ _6012_/A vssd1 vssd1 vccd1 vccd1 _6169_/A sky130_fd_sc_hd__clkbuf_2
X_8310_ _8552_/A _8552_/B vssd1 vssd1 vccd1 vccd1 _8310_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_8_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8241_ _8527_/A _8242_/B vssd1 vssd1 vccd1 vccd1 _8363_/A sky130_fd_sc_hd__nor2_2
X_5453_ _5453_/A _5453_/B vssd1 vssd1 vccd1 vccd1 _5454_/B sky130_fd_sc_hd__nand2_1
XFILLER_8_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4404_ _4407_/A vssd1 vssd1 vccd1 vccd1 _4404_/Y sky130_fd_sc_hd__inv_2
X_8172_ _8172_/A _8172_/B vssd1 vssd1 vccd1 vccd1 _8264_/A sky130_fd_sc_hd__nor2_2
X_5384_ _8695_/Q vssd1 vssd1 vccd1 vccd1 _6528_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_99_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7123_ _7123_/A _7123_/B _7123_/C vssd1 vssd1 vccd1 vccd1 _7139_/A sky130_fd_sc_hd__and3_1
X_7054_ _7231_/A _7225_/B vssd1 vssd1 vccd1 vccd1 _7056_/A sky130_fd_sc_hd__xnor2_1
X_6005_ _6274_/A _5986_/B _6180_/B vssd1 vssd1 vccd1 vccd1 _6323_/A sky130_fd_sc_hd__o21ai_4
XFILLER_55_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7956_ _8044_/B _7956_/B vssd1 vssd1 vccd1 vccd1 _7957_/B sky130_fd_sc_hd__nor2_1
X_7887_ _8139_/A _7887_/B vssd1 vssd1 vccd1 vccd1 _7887_/Y sky130_fd_sc_hd__nand2_1
X_6907_ _7020_/B _6873_/A _6873_/B _7400_/A _7118_/B vssd1 vssd1 vccd1 vccd1 _6907_/Y
+ sky130_fd_sc_hd__o32ai_2
XFILLER_35_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6838_ _6965_/A _6877_/A _6960_/B _6779_/B vssd1 vssd1 vccd1 vccd1 _6881_/A sky130_fd_sc_hd__a2bb2o_2
XFILLER_23_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8508_ _8445_/A _8444_/B _8442_/X vssd1 vssd1 vccd1 vccd1 _8509_/B sky130_fd_sc_hd__a21o_1
X_6769_ _6769_/A vssd1 vssd1 vccd1 vccd1 _7118_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_10_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8439_ _8439_/A _8531_/A _8439_/C vssd1 vssd1 vccd1 vccd1 _8443_/B sky130_fd_sc_hd__and3_1
XFILLER_104_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8795__12 vssd1 vssd1 vccd1 vccd1 _8795__12/HI _8890_/A sky130_fd_sc_hd__conb_1
X_7810_ _7813_/A _7813_/B _7813_/C vssd1 vssd1 vccd1 vccd1 _8381_/B sky130_fd_sc_hd__and3_1
XFILLER_91_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7741_ _8155_/A _7745_/A vssd1 vssd1 vccd1 vccd1 _7998_/A sky130_fd_sc_hd__nand2_2
X_4953_ _5215_/B _5142_/C _4953_/C vssd1 vssd1 vccd1 vccd1 _4953_/X sky130_fd_sc_hd__or3_1
X_7672_ _7672_/A _7672_/B vssd1 vssd1 vccd1 vccd1 _7762_/B sky130_fd_sc_hd__nand2_1
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6623_ _6798_/A vssd1 vssd1 vccd1 vccd1 _6793_/A sky130_fd_sc_hd__clkbuf_2
X_4884_ _4814_/D _4879_/X _5178_/B _4883_/Y vssd1 vssd1 vccd1 vccd1 _5291_/A sky130_fd_sc_hd__a211o_1
XFILLER_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6554_ _6583_/B vssd1 vssd1 vccd1 vccd1 _6588_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_5505_ _5505_/A _5505_/B vssd1 vssd1 vccd1 vccd1 _5530_/A sky130_fd_sc_hd__nand2_4
X_6485_ _6485_/A _6485_/B vssd1 vssd1 vccd1 vccd1 _8731_/D sky130_fd_sc_hd__nor2_1
X_8224_ _8229_/A _8229_/B vssd1 vssd1 vccd1 vccd1 _8225_/B sky130_fd_sc_hd__xor2_2
X_5436_ _5478_/A _5484_/A _5435_/X _8713_/Q vssd1 vssd1 vccd1 vccd1 _5436_/Y sky130_fd_sc_hd__a31oi_1
XFILLER_10_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8155_ _8155_/A _8155_/B _8155_/C vssd1 vssd1 vccd1 vccd1 _8173_/B sky130_fd_sc_hd__and3_1
X_5367_ _5372_/C _5367_/B _5389_/B vssd1 vssd1 vccd1 vccd1 _5368_/A sky130_fd_sc_hd__and3b_1
XFILLER_87_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8086_ _8086_/A _8086_/B vssd1 vssd1 vccd1 vccd1 _8147_/B sky130_fd_sc_hd__xor2_2
X_7106_ _7391_/A _7078_/A _7105_/Y vssd1 vssd1 vccd1 vccd1 _7126_/B sky130_fd_sc_hd__a21o_1
X_5298_ _5298_/A _5298_/B _5298_/C _5298_/D vssd1 vssd1 vccd1 vccd1 _5305_/C sky130_fd_sc_hd__or4_1
XFILLER_101_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7037_ _7037_/A _7200_/B vssd1 vssd1 vccd1 vccd1 _7038_/B sky130_fd_sc_hd__xnor2_1
XFILLER_74_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8988_ _8988_/A _4485_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[37] sky130_fd_sc_hd__ebufn_8
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7939_ _8102_/B vssd1 vssd1 vccd1 vccd1 _8098_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_82_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6270_ _6274_/A _6187_/B _6186_/A vssd1 vssd1 vccd1 vccd1 _6271_/B sky130_fd_sc_hd__a21oi_2
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5221_ _5221_/A _5221_/B _5221_/C _5220_/X vssd1 vssd1 vccd1 vccd1 _5221_/X sky130_fd_sc_hd__or4b_1
XFILLER_69_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5152_ _5259_/D _5151_/X _5271_/A vssd1 vssd1 vccd1 vccd1 _5152_/X sky130_fd_sc_hd__o21ba_1
XFILLER_69_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5083_ _5083_/A _5083_/B vssd1 vssd1 vccd1 vccd1 _5156_/B sky130_fd_sc_hd__nor2_2
X_8911_ _8911_/A _4394_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[30] sky130_fd_sc_hd__ebufn_8
XFILLER_49_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8773_ _8784_/CLK _8773_/D vssd1 vssd1 vccd1 vccd1 _8773_/Q sky130_fd_sc_hd__dfxtp_1
X_5985_ _5986_/B _6093_/A _5595_/Y vssd1 vssd1 vccd1 vccd1 _6185_/A sky130_fd_sc_hd__o21a_1
X_7724_ _8657_/Q _7734_/A vssd1 vssd1 vccd1 vccd1 _7725_/B sky130_fd_sc_hd__and2b_1
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4936_ _5215_/C _5263_/C vssd1 vssd1 vccd1 vccd1 _5108_/B sky130_fd_sc_hd__or2_2
X_7655_ _7654_/A _7654_/B _7654_/C vssd1 vssd1 vccd1 vccd1 _7656_/C sky130_fd_sc_hd__a21o_1
XFILLER_20_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4867_ _5083_/A _4867_/B vssd1 vssd1 vccd1 vccd1 _5048_/A sky130_fd_sc_hd__nor2_1
XFILLER_32_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6606_ _7589_/A _6606_/B _6606_/C vssd1 vssd1 vccd1 vccd1 _6607_/A sky130_fd_sc_hd__and3_1
X_7586_ _7579_/Y _7585_/X _7586_/S vssd1 vssd1 vccd1 vccd1 _7587_/C sky130_fd_sc_hd__mux2_1
XFILLER_20_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6537_ _7587_/A _6560_/A _7579_/B vssd1 vssd1 vccd1 vccd1 _6537_/X sky130_fd_sc_hd__o21a_1
X_4798_ _4798_/A vssd1 vssd1 vccd1 vccd1 _8667_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6468_ _8727_/Q _8726_/Q _8725_/Q vssd1 vssd1 vccd1 vccd1 _6473_/B sky130_fd_sc_hd__and3_1
X_8207_ _8232_/A _8207_/B vssd1 vssd1 vccd1 vccd1 _8223_/A sky130_fd_sc_hd__xnor2_2
X_6399_ _5709_/Y _6398_/B _6398_/Y _6390_/A _6390_/B vssd1 vssd1 vccd1 vccd1 _6399_/X
+ sky130_fd_sc_hd__a2111o_1
X_5419_ _8705_/Q vssd1 vssd1 vccd1 vccd1 _6415_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_87_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8138_ _8138_/A _8139_/B _8556_/A _8137_/X vssd1 vssd1 vccd1 vccd1 _8559_/B sky130_fd_sc_hd__or4bb_2
X_8069_ _8153_/B _8181_/A vssd1 vssd1 vccd1 vccd1 _8070_/B sky130_fd_sc_hd__xnor2_1
XFILLER_75_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5770_ _8713_/Q _7943_/B vssd1 vssd1 vccd1 vccd1 _5770_/Y sky130_fd_sc_hd__nor2_1
XFILLER_22_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4721_ _4995_/A vssd1 vssd1 vccd1 vccd1 _5271_/B sky130_fd_sc_hd__clkbuf_2
X_4652_ _8642_/Q _8641_/Q _4652_/C vssd1 vssd1 vccd1 vccd1 _4656_/B sky130_fd_sc_hd__and3_1
X_7440_ _7524_/S _7523_/A _7523_/B _7439_/Y vssd1 vssd1 vccd1 vccd1 _7514_/A sky130_fd_sc_hd__a31o_2
X_4583_ _4583_/A vssd1 vssd1 vccd1 vccd1 _8929_/A sky130_fd_sc_hd__clkbuf_1
X_7371_ _7335_/A _7335_/B _7370_/X vssd1 vssd1 vccd1 vccd1 _7483_/B sky130_fd_sc_hd__a21oi_2
X_6322_ _6275_/S _6276_/A _6321_/X vssd1 vssd1 vccd1 vccd1 _6325_/A sky130_fd_sc_hd__a21bo_1
Xclkbuf_4_5_0_wb_clk_i clkbuf_4_5_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _8723_/CLK
+ sky130_fd_sc_hd__clkbuf_2
X_6253_ _6337_/A _6253_/B vssd1 vssd1 vccd1 vccd1 _6255_/C sky130_fd_sc_hd__nor2_1
XFILLER_103_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5204_ _5197_/X _5203_/X _5224_/C vssd1 vssd1 vccd1 vccd1 _5204_/X sky130_fd_sc_hd__a21o_1
X_6184_ _6185_/B _6185_/C _6185_/A vssd1 vssd1 vccd1 vccd1 _6186_/A sky130_fd_sc_hd__o21a_1
XFILLER_69_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5135_ _5135_/A _5135_/B _5135_/C vssd1 vssd1 vccd1 vccd1 _5251_/C sky130_fd_sc_hd__or3_1
X_5066_ _5066_/A _5066_/B vssd1 vssd1 vccd1 vccd1 _5066_/Y sky130_fd_sc_hd__nand2_1
XFILLER_84_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5968_ _5957_/A _5957_/B _5967_/X vssd1 vssd1 vccd1 vccd1 _6129_/A sky130_fd_sc_hd__a21o_1
XFILLER_80_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8756_ _8758_/CLK _8756_/D vssd1 vssd1 vccd1 vccd1 _8756_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7707_ _8099_/A _7839_/B _7706_/Y vssd1 vssd1 vccd1 vccd1 _7711_/A sky130_fd_sc_hd__a21oi_1
X_4919_ _5190_/A _5004_/A vssd1 vssd1 vccd1 vccd1 _5098_/B sky130_fd_sc_hd__or2_1
X_5899_ _5837_/A _6183_/B _5838_/B _6004_/B vssd1 vssd1 vccd1 vccd1 _5903_/A sky130_fd_sc_hd__a2bb2o_1
X_8687_ _8704_/CLK _8687_/D vssd1 vssd1 vccd1 vccd1 _8687_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7638_ _7638_/A _7638_/B vssd1 vssd1 vccd1 vccd1 _7652_/C sky130_fd_sc_hd__nor2_1
XFILLER_20_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7569_ _7569_/A _7569_/B vssd1 vssd1 vccd1 vccd1 _7569_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_4_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6940_ _6940_/A _6940_/B vssd1 vssd1 vccd1 vccd1 _6996_/B sky130_fd_sc_hd__xor2_1
XFILLER_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6871_ _6871_/A _6870_/X vssd1 vssd1 vccd1 vccd1 _6875_/A sky130_fd_sc_hd__or2b_1
X_5822_ _5822_/A _5890_/B _5822_/C vssd1 vssd1 vccd1 vccd1 _5889_/A sky130_fd_sc_hd__nand3_1
X_8610_ _8782_/Q _8609_/A _8609_/Y _7642_/X vssd1 vssd1 vccd1 vccd1 _8782_/D sky130_fd_sc_hd__o211a_1
XFILLER_62_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8541_ _8236_/C _8356_/B _8358_/B vssd1 vssd1 vccd1 vccd1 _8542_/B sky130_fd_sc_hd__a21bo_1
X_5753_ _5754_/A _5754_/B _5754_/C vssd1 vssd1 vccd1 vccd1 _5845_/A sky130_fd_sc_hd__o21a_1
XFILLER_62_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4704_ _4747_/B vssd1 vssd1 vccd1 vccd1 _4760_/A sky130_fd_sc_hd__clkbuf_1
X_8472_ _8472_/A _8472_/B vssd1 vssd1 vccd1 vccd1 _8488_/B sky130_fd_sc_hd__xor2_1
X_5684_ _5684_/A _5684_/B vssd1 vssd1 vccd1 vccd1 _5684_/Y sky130_fd_sc_hd__nor2_1
X_7423_ _7423_/A _7423_/B vssd1 vssd1 vccd1 vccd1 _7425_/A sky130_fd_sc_hd__xnor2_1
X_4635_ _8636_/Q _4637_/C _4628_/X vssd1 vssd1 vccd1 vccd1 _4636_/B sky130_fd_sc_hd__o21ai_1
X_7354_ _7322_/B _7354_/B vssd1 vssd1 vccd1 vccd1 _7354_/X sky130_fd_sc_hd__and2b_1
X_4566_ _4566_/A _4566_/B _4695_/B vssd1 vssd1 vccd1 vccd1 _4574_/B sky130_fd_sc_hd__or3b_1
X_6305_ _6237_/A _6305_/B vssd1 vssd1 vccd1 vccd1 _6305_/X sky130_fd_sc_hd__and2b_1
XFILLER_103_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4497_ _8657_/Q vssd1 vssd1 vccd1 vccd1 _6615_/B sky130_fd_sc_hd__clkbuf_4
X_7285_ _7416_/A _7285_/B vssd1 vssd1 vccd1 vccd1 _7286_/B sky130_fd_sc_hd__nor2_1
X_6236_ _6154_/A _6154_/B _6235_/X vssd1 vssd1 vccd1 vccd1 _6305_/B sky130_fd_sc_hd__a21bo_1
X_6167_ _5921_/B _6173_/A _6166_/X vssd1 vssd1 vccd1 vccd1 _6168_/B sky130_fd_sc_hd__o21a_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5118_ _5188_/A _5118_/B vssd1 vssd1 vccd1 vccd1 _5190_/C sky130_fd_sc_hd__nand2_1
X_6098_ _6099_/A _6099_/B vssd1 vssd1 vccd1 vccd1 _6207_/B sky130_fd_sc_hd__or2_2
XFILLER_84_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5049_ _5135_/A _5136_/B vssd1 vssd1 vccd1 vccd1 _5126_/D sky130_fd_sc_hd__or2_1
XFILLER_72_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8739_ _8742_/CLK _8739_/D vssd1 vssd1 vccd1 vccd1 _8739_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4420_ _4426_/A vssd1 vssd1 vccd1 vccd1 _4425_/A sky130_fd_sc_hd__buf_4
XFILLER_8_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7070_ _7070_/A _7070_/B vssd1 vssd1 vccd1 vccd1 _7086_/B sky130_fd_sc_hd__xnor2_1
XFILLER_100_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6021_ _6250_/A vssd1 vssd1 vccd1 vccd1 _6058_/A sky130_fd_sc_hd__inv_2
XFILLER_86_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7972_ _7972_/A _7972_/B _7972_/C vssd1 vssd1 vccd1 vccd1 _7974_/A sky130_fd_sc_hd__nor3_1
XFILLER_54_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6923_ _7034_/A vssd1 vssd1 vccd1 vccd1 _7391_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_22_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6854_ _6854_/A vssd1 vssd1 vccd1 vccd1 _7182_/A sky130_fd_sc_hd__buf_2
XFILLER_35_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5805_ _5805_/A _5805_/B vssd1 vssd1 vccd1 vccd1 _5959_/A sky130_fd_sc_hd__nand2_1
XFILLER_13_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6785_ _6786_/A _6786_/B vssd1 vssd1 vccd1 vccd1 _6801_/B sky130_fd_sc_hd__nand2_1
X_8524_ _8461_/S _8460_/A _7999_/X vssd1 vssd1 vccd1 vccd1 _8525_/B sky130_fd_sc_hd__a21oi_1
X_5736_ _5634_/A _5735_/X _5634_/C _5619_/A vssd1 vssd1 vccd1 vccd1 _5983_/A sky130_fd_sc_hd__a31o_1
X_8455_ _8371_/A _8371_/B _8370_/A vssd1 vssd1 vccd1 vccd1 _8456_/B sky130_fd_sc_hd__a21oi_2
X_5667_ _5667_/A _5667_/B vssd1 vssd1 vccd1 vccd1 _5670_/A sky130_fd_sc_hd__xnor2_1
X_4618_ _4640_/A vssd1 vssd1 vccd1 vccd1 _4679_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7406_ _7406_/A _7284_/A vssd1 vssd1 vccd1 vccd1 _7406_/X sky130_fd_sc_hd__or2b_1
X_8386_ _8386_/A _8386_/B vssd1 vssd1 vccd1 vccd1 _8387_/C sky130_fd_sc_hd__nand2_1
X_5598_ _5678_/A _5678_/B vssd1 vssd1 vccd1 vccd1 _5679_/A sky130_fd_sc_hd__or2_1
XFILLER_89_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7337_ _7235_/A _7235_/B _7336_/Y vssd1 vssd1 vccd1 vccd1 _7338_/B sky130_fd_sc_hd__o21a_1
XFILLER_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4549_ _4549_/A _4814_/C _4574_/A _4568_/C vssd1 vssd1 vccd1 vccd1 _4550_/A sky130_fd_sc_hd__or4_4
XFILLER_104_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7268_ _7268_/A _7268_/B _7268_/C vssd1 vssd1 vccd1 vccd1 _7409_/A sky130_fd_sc_hd__nand3_1
XFILLER_104_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6219_ _6161_/A _6219_/B vssd1 vssd1 vccd1 vccd1 _6219_/X sky130_fd_sc_hd__and2b_1
XFILLER_89_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_10 _4947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7199_ _7023_/A _7023_/B _7198_/X vssd1 vssd1 vccd1 vccd1 _7325_/B sky130_fd_sc_hd__a21bo_1
XFILLER_38_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6570_ _6570_/A _8747_/Q vssd1 vssd1 vccd1 vccd1 _6572_/B sky130_fd_sc_hd__xor2_1
X_5521_ _5521_/A _5521_/B vssd1 vssd1 vccd1 vccd1 _6012_/A sky130_fd_sc_hd__xnor2_2
X_8240_ _8496_/S _8239_/X _8192_/Y vssd1 vssd1 vccd1 vccd1 _8242_/B sky130_fd_sc_hd__a21o_1
XFILLER_8_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5452_ _5452_/A _8706_/Q vssd1 vssd1 vccd1 vccd1 _5453_/B sky130_fd_sc_hd__or2b_1
XFILLER_99_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4403_ _4407_/A vssd1 vssd1 vccd1 vccd1 _4403_/Y sky130_fd_sc_hd__inv_2
X_8171_ _8450_/A _8248_/B vssd1 vssd1 vccd1 vccd1 _8175_/A sky130_fd_sc_hd__nand2_1
X_5383_ _5387_/C _5383_/B vssd1 vssd1 vccd1 vccd1 _8694_/D sky130_fd_sc_hd__nor2_1
X_7122_ _7134_/A _7122_/B vssd1 vssd1 vccd1 vccd1 _7140_/B sky130_fd_sc_hd__nor2_1
XFILLER_101_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7053_ _7227_/A _7227_/B vssd1 vssd1 vccd1 vccd1 _7225_/B sky130_fd_sc_hd__xnor2_1
XFILLER_5_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6004_ _6004_/A _6004_/B vssd1 vssd1 vccd1 vccd1 _6180_/B sky130_fd_sc_hd__nand2_2
XFILLER_67_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7955_ _7955_/A _7955_/B vssd1 vssd1 vccd1 vccd1 _7956_/B sky130_fd_sc_hd__and2_1
XFILLER_42_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7886_ _8586_/A _7889_/A vssd1 vssd1 vccd1 vccd1 _7887_/B sky130_fd_sc_hd__nand2_1
X_6906_ _7279_/B vssd1 vssd1 vccd1 vccd1 _7400_/A sky130_fd_sc_hd__buf_2
XFILLER_50_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6837_ _7118_/A _6837_/B vssd1 vssd1 vccd1 vccd1 _6877_/A sky130_fd_sc_hd__nand2_1
X_8507_ _8433_/A _8433_/B _8506_/X vssd1 vssd1 vccd1 vccd1 _8510_/A sky130_fd_sc_hd__a21oi_2
X_6768_ _6768_/A vssd1 vssd1 vccd1 vccd1 _6769_/A sky130_fd_sc_hd__inv_2
X_5719_ _5984_/C vssd1 vssd1 vccd1 vccd1 _5986_/A sky130_fd_sc_hd__inv_2
X_6699_ _7392_/B vssd1 vssd1 vccd1 vccd1 _6949_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_40_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8438_ _8372_/B _8438_/B vssd1 vssd1 vccd1 vccd1 _8443_/A sky130_fd_sc_hd__and2b_1
X_8369_ _8369_/A _8369_/B vssd1 vssd1 vccd1 vccd1 _8370_/B sky130_fd_sc_hd__nor2_1
XFILLER_2_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7740_ _7821_/A _7821_/B vssd1 vssd1 vccd1 vccd1 _7745_/A sky130_fd_sc_hd__nand2_2
XFILLER_51_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4952_ _5215_/C vssd1 vssd1 vccd1 vccd1 _5142_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_36_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7671_ _7671_/A vssd1 vssd1 vccd1 vccd1 _7762_/A sky130_fd_sc_hd__buf_2
X_4883_ _4883_/A _4883_/B vssd1 vssd1 vccd1 vccd1 _4883_/Y sky130_fd_sc_hd__nor2_1
X_6622_ _6645_/A _6645_/B vssd1 vssd1 vccd1 vccd1 _6798_/A sky130_fd_sc_hd__and2_1
X_6553_ _8747_/Q vssd1 vssd1 vccd1 vccd1 _6583_/B sky130_fd_sc_hd__inv_2
X_5504_ _5493_/A _5526_/B _5500_/X _5498_/X vssd1 vssd1 vccd1 vccd1 _5505_/B sky130_fd_sc_hd__a211o_1
X_6484_ _6482_/A _6486_/C _6483_/X vssd1 vssd1 vccd1 vccd1 _6485_/B sky130_fd_sc_hd__o21ai_1
X_8223_ _8223_/A _8223_/B vssd1 vssd1 vccd1 vccd1 _8229_/B sky130_fd_sc_hd__xnor2_2
X_5435_ _5452_/A _8707_/Q _5463_/B _5456_/B vssd1 vssd1 vccd1 vccd1 _5435_/X sky130_fd_sc_hd__a211o_1
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8154_ _8371_/A _8070_/B _8153_/X vssd1 vssd1 vccd1 vccd1 _8256_/A sky130_fd_sc_hd__a21o_1
X_5366_ _8687_/Q _6532_/B _5359_/B _8689_/Q vssd1 vssd1 vccd1 vccd1 _5367_/B sky130_fd_sc_hd__a31o_1
XFILLER_101_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8085_ _8182_/B _8082_/Y _8201_/A vssd1 vssd1 vccd1 vccd1 _8086_/B sky130_fd_sc_hd__a21oi_2
X_7105_ _7105_/A _7105_/B vssd1 vssd1 vccd1 vccd1 _7105_/Y sky130_fd_sc_hd__nor2_1
X_5297_ _4541_/X _4549_/A _4925_/A vssd1 vssd1 vccd1 vccd1 _5298_/D sky130_fd_sc_hd__o21a_1
X_7036_ _7036_/A _7331_/A vssd1 vssd1 vccd1 vccd1 _7200_/B sky130_fd_sc_hd__xnor2_1
XFILLER_19_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8987_ _8987_/A _4484_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[36] sky130_fd_sc_hd__ebufn_8
XFILLER_82_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7938_ _7938_/A _7938_/B vssd1 vssd1 vccd1 vccd1 _8036_/A sky130_fd_sc_hd__nor2_1
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7869_ _7976_/A _7869_/B vssd1 vssd1 vccd1 vccd1 _7891_/B sky130_fd_sc_hd__nand2_1
XFILLER_50_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5220_ _5207_/Y _5210_/B _5280_/A vssd1 vssd1 vccd1 vccd1 _5220_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8855__72 vssd1 vssd1 vccd1 vccd1 _8855__72/HI _8964_/A sky130_fd_sc_hd__conb_1
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5151_ _4823_/A _5145_/Y _5148_/X _5150_/A _5150_/Y vssd1 vssd1 vccd1 vccd1 _5151_/X
+ sky130_fd_sc_hd__a221o_1
X_5082_ _5083_/A _5082_/B vssd1 vssd1 vccd1 vccd1 _5188_/B sky130_fd_sc_hd__nor2_2
X_8910_ _8910_/A _4393_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[29] sky130_fd_sc_hd__ebufn_8
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8772_ _8784_/CLK _8772_/D vssd1 vssd1 vccd1 vccd1 _8772_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5984_ _6192_/B _6262_/B _5984_/C vssd1 vssd1 vccd1 vccd1 _6093_/A sky130_fd_sc_hd__and3b_1
X_7723_ _8781_/Q _8657_/Q vssd1 vssd1 vccd1 vccd1 _7725_/A sky130_fd_sc_hd__and2b_1
XFILLER_52_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4935_ _4935_/A _4935_/B vssd1 vssd1 vccd1 vccd1 _5263_/C sky130_fd_sc_hd__nor2_2
XFILLER_60_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7654_ _7654_/A _7654_/B _7654_/C vssd1 vssd1 vccd1 vccd1 _7666_/S sky130_fd_sc_hd__and3_1
XFILLER_20_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4866_ _4541_/X _4897_/C _4901_/B _5083_/B vssd1 vssd1 vccd1 vccd1 _4867_/B sky130_fd_sc_hd__o31a_1
X_7585_ _7585_/A _7585_/B vssd1 vssd1 vccd1 vccd1 _7585_/X sky130_fd_sc_hd__or2_1
X_4797_ _4804_/C _7576_/B _4797_/C vssd1 vssd1 vccd1 vccd1 _4798_/A sky130_fd_sc_hd__and3b_1
X_6605_ _7583_/B _6604_/C _6851_/A vssd1 vssd1 vccd1 vccd1 _6606_/C sky130_fd_sc_hd__o21ai_1
XFILLER_21_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6536_ _8746_/Q vssd1 vssd1 vccd1 vccd1 _7579_/B sky130_fd_sc_hd__clkbuf_2
X_6467_ _8726_/Q _6455_/B _6466_/Y vssd1 vssd1 vccd1 vccd1 _8726_/D sky130_fd_sc_hd__o21a_1
X_8206_ _8206_/A _8206_/B vssd1 vssd1 vccd1 vccd1 _8207_/B sky130_fd_sc_hd__xor2_2
X_6398_ _6398_/A _6398_/B vssd1 vssd1 vccd1 vccd1 _6398_/Y sky130_fd_sc_hd__nor2_1
X_5418_ _8721_/Q vssd1 vssd1 vccd1 vccd1 _6415_/A sky130_fd_sc_hd__inv_2
XFILLER_102_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8137_ _8053_/B _8053_/C _8053_/A vssd1 vssd1 vccd1 vccd1 _8137_/X sky130_fd_sc_hd__a21o_1
X_5349_ _8684_/Q _5349_/B vssd1 vssd1 vccd1 vccd1 _8684_/D sky130_fd_sc_hd__nor2_1
XFILLER_101_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8068_ _8068_/A _8068_/B vssd1 vssd1 vccd1 vccd1 _8181_/A sky130_fd_sc_hd__xnor2_2
XFILLER_101_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7019_ _7019_/A _7185_/A vssd1 vssd1 vccd1 vccd1 _7417_/A sky130_fd_sc_hd__xnor2_4
XFILLER_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4720_ _4720_/A vssd1 vssd1 vccd1 vccd1 _4995_/A sky130_fd_sc_hd__clkbuf_2
X_4651_ _8641_/Q _4652_/C _4650_/Y vssd1 vssd1 vccd1 vccd1 _8641_/D sky130_fd_sc_hd__a21oi_1
X_4582_ _8675_/Q _4584_/B vssd1 vssd1 vccd1 vccd1 _4583_/A sky130_fd_sc_hd__and2_1
X_7370_ _7370_/A _7370_/B _7370_/C vssd1 vssd1 vccd1 vccd1 _7370_/X sky130_fd_sc_hd__and3_1
X_6321_ _6263_/A _5897_/A _6275_/S _6276_/A _6276_/B vssd1 vssd1 vccd1 vccd1 _6321_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_89_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6252_ _6252_/A _6252_/B _6311_/B vssd1 vssd1 vccd1 vccd1 _6253_/B sky130_fd_sc_hd__and3_1
X_6183_ _6183_/A _6183_/B vssd1 vssd1 vccd1 vccd1 _6185_/B sky130_fd_sc_hd__nor2_1
X_5203_ _5059_/B _5219_/A _5200_/X _5202_/X _4702_/D vssd1 vssd1 vccd1 vccd1 _5203_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_69_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5134_ _5154_/A vssd1 vssd1 vccd1 vccd1 _5250_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_84_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5065_ _5176_/A _5272_/B _5056_/X _5064_/X _4818_/B vssd1 vssd1 vccd1 vccd1 _5073_/B
+ sky130_fd_sc_hd__o311a_1
XFILLER_84_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5967_ _5956_/B _5967_/B vssd1 vssd1 vccd1 vccd1 _5967_/X sky130_fd_sc_hd__and2b_1
XFILLER_80_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8755_ _8758_/CLK _8755_/D vssd1 vssd1 vccd1 vccd1 _8755_/Q sky130_fd_sc_hd__dfxtp_1
X_7706_ _7946_/A _8293_/A vssd1 vssd1 vccd1 vccd1 _7706_/Y sky130_fd_sc_hd__nor2_1
X_4918_ _5281_/B _5183_/A vssd1 vssd1 vccd1 vccd1 _5004_/A sky130_fd_sc_hd__or2_1
X_8686_ _8704_/CLK _8686_/D vssd1 vssd1 vccd1 vccd1 _8686_/Q sky130_fd_sc_hd__dfxtp_1
X_5898_ _5975_/A _5975_/B vssd1 vssd1 vccd1 vccd1 _5905_/A sky130_fd_sc_hd__xnor2_1
X_7637_ _7637_/A _7637_/B vssd1 vssd1 vccd1 vccd1 _7638_/B sky130_fd_sc_hd__and2_1
X_4849_ _4877_/B _4872_/B vssd1 vssd1 vccd1 vccd1 _4901_/B sky130_fd_sc_hd__nand2_1
X_7568_ _7565_/A _7565_/B _7563_/A vssd1 vssd1 vccd1 vccd1 _7569_/B sky130_fd_sc_hd__a21oi_1
X_7499_ _7499_/A _7499_/B vssd1 vssd1 vccd1 vccd1 _7500_/B sky130_fd_sc_hd__xnor2_1
X_6519_ _8743_/Q _6519_/B vssd1 vssd1 vccd1 vccd1 _6521_/A sky130_fd_sc_hd__and2_1
XFILLER_0_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8825__42 vssd1 vssd1 vccd1 vccd1 _8825__42/HI _8920_/A sky130_fd_sc_hd__conb_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6870_ _6869_/B _6869_/C _6883_/A vssd1 vssd1 vccd1 vccd1 _6870_/X sky130_fd_sc_hd__a21o_1
X_5821_ _5820_/B _5890_/A _5986_/B vssd1 vssd1 vccd1 vccd1 _5822_/C sky130_fd_sc_hd__a21o_1
X_8540_ _8475_/A _8475_/B _8539_/Y vssd1 vssd1 vccd1 vccd1 _8542_/A sky130_fd_sc_hd__o21ai_1
X_5752_ _5835_/A _6004_/B vssd1 vssd1 vccd1 vccd1 _5754_/C sky130_fd_sc_hd__xnor2_1
X_4703_ _6460_/A _4771_/B vssd1 vssd1 vccd1 vccd1 _4747_/B sky130_fd_sc_hd__and2_1
X_8471_ _8471_/A _8471_/B vssd1 vssd1 vccd1 vccd1 _8472_/B sky130_fd_sc_hd__xnor2_2
X_5683_ _5683_/A _5683_/B vssd1 vssd1 vccd1 vccd1 _5684_/B sky130_fd_sc_hd__and2_1
XFILLER_30_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7422_ _7487_/A _7487_/B vssd1 vssd1 vccd1 vccd1 _7423_/B sky130_fd_sc_hd__xor2_1
X_4634_ _8636_/Q _4637_/C vssd1 vssd1 vccd1 vccd1 _4636_/A sky130_fd_sc_hd__and2_1
X_4565_ _5249_/A _4565_/B vssd1 vssd1 vccd1 vccd1 _4695_/B sky130_fd_sc_hd__nor2_1
X_7353_ _7340_/A _7340_/B _7352_/X vssd1 vssd1 vccd1 vccd1 _7432_/A sky130_fd_sc_hd__a21bo_2
X_6304_ _6304_/A _6304_/B vssd1 vssd1 vccd1 vccd1 _6356_/A sky130_fd_sc_hd__xnor2_1
X_7284_ _7284_/A _7406_/A vssd1 vssd1 vccd1 vccd1 _7420_/A sky130_fd_sc_hd__xnor2_1
X_4496_ _6660_/B vssd1 vssd1 vccd1 vccd1 _5249_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6235_ _6235_/A _6155_/A vssd1 vssd1 vccd1 vccd1 _6235_/X sky130_fd_sc_hd__or2b_1
XFILLER_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6166_ _6166_/A _6312_/S vssd1 vssd1 vccd1 vccd1 _6166_/X sky130_fd_sc_hd__or2_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6097_ _6190_/A _6190_/B vssd1 vssd1 vccd1 vccd1 _6099_/B sky130_fd_sc_hd__xnor2_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5117_ _5108_/B _5117_/B vssd1 vssd1 vccd1 vccd1 _5118_/B sky130_fd_sc_hd__and2b_1
X_5048_ _5048_/A vssd1 vssd1 vccd1 vccd1 _5135_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_84_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6999_ _6999_/A _6905_/B vssd1 vssd1 vccd1 vccd1 _7000_/A sky130_fd_sc_hd__or2b_1
X_8738_ _8742_/CLK _8738_/D vssd1 vssd1 vccd1 vccd1 _8738_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8669_ _8771_/CLK _8669_/D vssd1 vssd1 vccd1 vccd1 _8669_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_5_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6020_ _5766_/A _5700_/C _5928_/B vssd1 vssd1 vccd1 vccd1 _6250_/A sky130_fd_sc_hd__o21ba_1
XFILLER_67_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7971_ _8051_/A _7971_/B vssd1 vssd1 vccd1 vccd1 _7972_/C sky130_fd_sc_hd__nand2_1
XFILLER_81_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6922_ _6922_/A _6922_/B vssd1 vssd1 vccd1 vccd1 _6938_/A sky130_fd_sc_hd__nand2_1
XFILLER_62_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6853_ _7036_/A _6646_/A _7011_/A vssd1 vssd1 vccd1 vccd1 _6854_/A sky130_fd_sc_hd__mux2_1
X_5804_ _5809_/B _5804_/B vssd1 vssd1 vccd1 vccd1 _5962_/B sky130_fd_sc_hd__xor2_2
XFILLER_35_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6784_ _6960_/B _6784_/B vssd1 vssd1 vccd1 vccd1 _6786_/B sky130_fd_sc_hd__xnor2_1
X_8523_ _7813_/A _7813_/C _7807_/B vssd1 vssd1 vccd1 vccd1 _8525_/A sky130_fd_sc_hd__a21o_1
X_5735_ _6433_/A _6653_/B vssd1 vssd1 vccd1 vccd1 _5735_/X sky130_fd_sc_hd__or2_1
XFILLER_50_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8454_ _8528_/A _8528_/B vssd1 vssd1 vccd1 vccd1 _8456_/A sky130_fd_sc_hd__xnor2_2
X_5666_ _5666_/A _5666_/B vssd1 vssd1 vccd1 vccd1 _5667_/B sky130_fd_sc_hd__xnor2_1
X_4617_ _5462_/A input2/X vssd1 vssd1 vccd1 vccd1 _4640_/A sky130_fd_sc_hd__and2b_1
X_7405_ _7405_/A _7497_/A vssd1 vssd1 vccd1 vccd1 _7457_/B sky130_fd_sc_hd__xnor2_1
X_8385_ _8459_/B _8384_/C _8384_/A vssd1 vssd1 vccd1 vccd1 _8387_/B sky130_fd_sc_hd__a21o_1
X_5597_ _5749_/A _5597_/B vssd1 vssd1 vccd1 vccd1 _5678_/B sky130_fd_sc_hd__xnor2_1
X_7336_ _7336_/A _7336_/B vssd1 vssd1 vccd1 vccd1 _7336_/Y sky130_fd_sc_hd__nand2_1
X_4548_ _7943_/B _4814_/B vssd1 vssd1 vccd1 vccd1 _4568_/C sky130_fd_sc_hd__nand2_1
XFILLER_104_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4479_ _4480_/A vssd1 vssd1 vccd1 vccd1 _4479_/Y sky130_fd_sc_hd__inv_2
X_7267_ _7266_/B _7266_/C _7280_/S vssd1 vssd1 vccd1 vccd1 _7268_/C sky130_fd_sc_hd__a21o_1
X_6218_ _6215_/A _6218_/B vssd1 vssd1 vccd1 vccd1 _6290_/B sky130_fd_sc_hd__and2b_1
X_7198_ _7198_/A _7198_/B _7198_/C vssd1 vssd1 vccd1 vccd1 _7198_/X sky130_fd_sc_hd__or3_1
XFILLER_97_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6149_ _5920_/A _6227_/A _6149_/C vssd1 vssd1 vccd1 vccd1 _6227_/B sky130_fd_sc_hd__nand3b_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_11 _5088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5520_ _5518_/X _5544_/A vssd1 vssd1 vccd1 vccd1 _5521_/B sky130_fd_sc_hd__and2b_1
X_5451_ _8706_/Q _5452_/A vssd1 vssd1 vccd1 vccd1 _5453_/A sky130_fd_sc_hd__or2b_1
X_4402_ _4426_/A vssd1 vssd1 vccd1 vccd1 _4407_/A sky130_fd_sc_hd__buf_6
X_8170_ _8256_/A _8256_/B vssd1 vssd1 vccd1 vccd1 _8179_/A sky130_fd_sc_hd__xnor2_2
X_5382_ _8694_/Q _5381_/B _5360_/X vssd1 vssd1 vccd1 vccd1 _5383_/B sky130_fd_sc_hd__o21ai_1
X_7121_ _6825_/A _7120_/B _6809_/A vssd1 vssd1 vccd1 vccd1 _7122_/B sky130_fd_sc_hd__o21a_1
XFILLER_101_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7052_ _7331_/A _7052_/B vssd1 vssd1 vccd1 vccd1 _7227_/B sky130_fd_sc_hd__xnor2_1
X_6003_ _6004_/B vssd1 vssd1 vccd1 vccd1 _6274_/A sky130_fd_sc_hd__buf_2
XFILLER_27_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7954_ _7955_/A _7955_/B vssd1 vssd1 vccd1 vccd1 _8044_/B sky130_fd_sc_hd__nor2_1
XFILLER_27_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6905_ _6999_/A _6905_/B vssd1 vssd1 vccd1 vccd1 _6918_/A sky130_fd_sc_hd__xnor2_1
X_7885_ _8586_/A _7889_/A vssd1 vssd1 vccd1 vccd1 _8139_/A sky130_fd_sc_hd__or2_1
XFILLER_23_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6836_ _6836_/A _6910_/A vssd1 vssd1 vccd1 vccd1 _6837_/B sky130_fd_sc_hd__and2_1
X_6767_ _6786_/A _7119_/A _6767_/C vssd1 vssd1 vccd1 vccd1 _6963_/A sky130_fd_sc_hd__and3_1
X_8506_ _8429_/B _8506_/B vssd1 vssd1 vccd1 vccd1 _8506_/X sky130_fd_sc_hd__and2b_1
X_5718_ _5640_/A _5640_/B _5717_/X vssd1 vssd1 vccd1 vccd1 _5811_/A sky130_fd_sc_hd__a21o_1
XFILLER_10_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6698_ _7205_/B vssd1 vssd1 vccd1 vccd1 _7392_/B sky130_fd_sc_hd__clkbuf_2
X_8437_ _8527_/A _8437_/B vssd1 vssd1 vccd1 vccd1 _8445_/A sky130_fd_sc_hd__nor2_1
X_5649_ _8713_/Q _7842_/B vssd1 vssd1 vccd1 vccd1 _5650_/B sky130_fd_sc_hd__nand2_1
XFILLER_40_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8368_ _8369_/A _8369_/B vssd1 vssd1 vccd1 vccd1 _8370_/A sky130_fd_sc_hd__and2_1
XFILLER_104_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7319_ _7319_/A _7319_/B vssd1 vssd1 vccd1 vccd1 _7320_/B sky130_fd_sc_hd__nor2_1
XFILLER_104_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8299_ _8299_/A _8299_/B vssd1 vssd1 vccd1 vccd1 _8300_/B sky130_fd_sc_hd__nand2_1
XFILLER_49_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4951_ _5077_/C vssd1 vssd1 vccd1 vccd1 _5215_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_36_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4882_ _5298_/C _4882_/B vssd1 vssd1 vccd1 vccd1 _5178_/B sky130_fd_sc_hd__nor2_1
X_7670_ _8665_/Q _8768_/Q vssd1 vssd1 vccd1 vccd1 _7671_/A sky130_fd_sc_hd__or2b_1
X_6621_ _6621_/A _6621_/B vssd1 vssd1 vccd1 vccd1 _6645_/B sky130_fd_sc_hd__nand2_1
X_6552_ _6628_/B _6570_/A _6583_/A vssd1 vssd1 vccd1 vccd1 _6552_/X sky130_fd_sc_hd__o21a_1
X_5503_ _5547_/A _5547_/B vssd1 vssd1 vccd1 vccd1 _5698_/A sky130_fd_sc_hd__xor2_2
X_6483_ _6508_/B vssd1 vssd1 vccd1 vccd1 _6483_/X sky130_fd_sc_hd__buf_2
X_8222_ _8222_/A _8222_/B vssd1 vssd1 vccd1 vccd1 _8223_/B sky130_fd_sc_hd__xor2_2
X_5434_ _8709_/Q vssd1 vssd1 vccd1 vccd1 _5456_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_8153_ _8181_/A _8153_/B vssd1 vssd1 vccd1 vccd1 _8153_/X sky130_fd_sc_hd__and2b_1
XFILLER_99_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5365_ _8689_/Q _8688_/Q _5365_/C vssd1 vssd1 vccd1 vccd1 _5372_/C sky130_fd_sc_hd__and3_1
X_7104_ _7104_/A _7104_/B vssd1 vssd1 vccd1 vccd1 _7126_/A sky130_fd_sc_hd__xor2_1
XFILLER_99_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8084_ _8082_/Y _8083_/X _8182_/B vssd1 vssd1 vccd1 vccd1 _8201_/A sky130_fd_sc_hd__a21oi_2
X_5296_ _5296_/A _5301_/C _5296_/C _5296_/D vssd1 vssd1 vccd1 vccd1 _5305_/B sky130_fd_sc_hd__or4_1
XFILLER_59_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7035_ _7035_/A vssd1 vssd1 vccd1 vccd1 _7331_/A sky130_fd_sc_hd__buf_2
XFILLER_19_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8986_ _8986_/A _4483_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[35] sky130_fd_sc_hd__ebufn_8
XFILLER_27_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7937_ _7981_/B _7981_/C _7981_/A vssd1 vssd1 vccd1 vccd1 _7964_/B sky130_fd_sc_hd__a21o_1
XFILLER_27_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7868_ _7893_/A _7867_/C _7867_/A vssd1 vssd1 vccd1 vccd1 _7869_/B sky130_fd_sc_hd__o21ai_1
Xclkbuf_2_0_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
X_6819_ _6820_/A _6820_/B vssd1 vssd1 vccd1 vccd1 _6953_/A sky130_fd_sc_hd__nor2_1
XFILLER_50_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7799_ _7799_/A _7799_/B vssd1 vssd1 vccd1 vccd1 _8273_/A sky130_fd_sc_hd__xnor2_2
XFILLER_7_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5150_ _5150_/A _5150_/B vssd1 vssd1 vccd1 vccd1 _5150_/Y sky130_fd_sc_hd__nor2_1
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5081_ _5159_/B _5149_/D vssd1 vssd1 vccd1 vccd1 _5228_/C sky130_fd_sc_hd__or2_1
X_8870__87 vssd1 vssd1 vccd1 vccd1 _8870__87/HI _8979_/A sky130_fd_sc_hd__conb_1
XFILLER_96_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5983_ _5983_/A vssd1 vssd1 vccd1 vccd1 _6192_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_64_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8771_ _8771_/CLK _8771_/D vssd1 vssd1 vccd1 vccd1 _8771_/Q sky130_fd_sc_hd__dfxtp_1
X_7722_ _7722_/A _7722_/B vssd1 vssd1 vccd1 vccd1 _7799_/A sky130_fd_sc_hd__nor2_4
X_4934_ _4934_/A _4934_/B vssd1 vssd1 vccd1 vccd1 _5215_/C sky130_fd_sc_hd__nor2_2
X_7653_ _7649_/A _7637_/B _7638_/B _7652_/X vssd1 vssd1 vccd1 vccd1 _7654_/C sky130_fd_sc_hd__a211o_1
X_4865_ _4901_/A _4897_/B _4897_/C _4778_/A vssd1 vssd1 vccd1 vccd1 _5083_/B sky130_fd_sc_hd__or4bb_2
X_4796_ _5501_/B _4796_/B vssd1 vssd1 vccd1 vccd1 _4797_/C sky130_fd_sc_hd__nand2_1
X_6604_ _6851_/A _7587_/B _6604_/C vssd1 vssd1 vccd1 vccd1 _6606_/B sky130_fd_sc_hd__or3_1
X_7584_ _7581_/Y _7582_/X _7583_/Y _5491_/X vssd1 vssd1 vccd1 vccd1 _8764_/D sky130_fd_sc_hd__o211ai_1
XFILLER_21_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6535_ _6535_/A _6535_/B _6535_/C _6535_/D vssd1 vssd1 vccd1 vccd1 _6560_/A sky130_fd_sc_hd__or4_4
X_8205_ _8302_/B _8205_/B vssd1 vssd1 vccd1 vccd1 _8206_/B sky130_fd_sc_hd__nor2_1
X_6466_ _8726_/Q _6455_/B _6465_/X vssd1 vssd1 vccd1 vccd1 _6466_/Y sky130_fd_sc_hd__a21boi_1
X_6397_ _6387_/X _6383_/X _6395_/X _6396_/Y vssd1 vssd1 vccd1 vccd1 _8716_/D sky130_fd_sc_hd__a31oi_1
X_5417_ _6409_/A _6405_/A _8721_/Q vssd1 vssd1 vccd1 vccd1 _5417_/X sky130_fd_sc_hd__o21a_1
X_8136_ _8311_/A _8311_/B vssd1 vssd1 vccd1 vccd1 _8556_/B sky130_fd_sc_hd__xor2_2
X_5348_ _6567_/A vssd1 vssd1 vccd1 vccd1 _5349_/B sky130_fd_sc_hd__inv_2
XFILLER_99_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8067_ _8380_/A _8064_/Y _8066_/X vssd1 vssd1 vccd1 vccd1 _8068_/B sky130_fd_sc_hd__a21boi_1
X_7018_ _6909_/S _6907_/Y _7017_/X vssd1 vssd1 vccd1 vccd1 _7023_/A sky130_fd_sc_hd__a21o_1
X_5279_ _5150_/A _5192_/B _5274_/X _5278_/X vssd1 vssd1 vccd1 vccd1 _5279_/X sky130_fd_sc_hd__o31a_1
XFILLER_28_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8969_ _8969_/A _4462_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[18] sky130_fd_sc_hd__ebufn_8
XFILLER_15_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4650_ _8641_/Q _4652_/C _4640_/X vssd1 vssd1 vccd1 vccd1 _4650_/Y sky130_fd_sc_hd__o21ai_1
X_4581_ _4581_/A vssd1 vssd1 vccd1 vccd1 _8928_/A sky130_fd_sc_hd__clkbuf_1
X_6320_ _6320_/A _6320_/B vssd1 vssd1 vccd1 vccd1 _6340_/A sky130_fd_sc_hd__xnor2_1
X_6251_ _6251_/A _6251_/B vssd1 vssd1 vccd1 vccd1 _6311_/B sky130_fd_sc_hd__nand2_1
XFILLER_97_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6182_ _6087_/A _6087_/B _6181_/Y vssd1 vssd1 vccd1 vccd1 _6188_/A sky130_fd_sc_hd__o21ai_2
X_5202_ _5202_/A _5227_/B vssd1 vssd1 vccd1 vccd1 _5202_/X sky130_fd_sc_hd__or2_1
XFILLER_69_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5133_ _4975_/X _4977_/Y _4997_/X _5132_/X vssd1 vssd1 vccd1 vccd1 _5133_/Y sky130_fd_sc_hd__o31ai_1
XFILLER_96_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5064_ _5192_/A _5250_/B _5064_/C _5071_/C vssd1 vssd1 vccd1 vccd1 _5064_/X sky130_fd_sc_hd__or4_1
XFILLER_37_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5966_ _6370_/A _5965_/Y _6370_/B vssd1 vssd1 vccd1 vccd1 _6367_/C sky130_fd_sc_hd__o21ai_1
XFILLER_13_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8754_ _8765_/CLK _8754_/D vssd1 vssd1 vccd1 vccd1 _8754_/Q sky130_fd_sc_hd__dfxtp_1
X_7705_ _7854_/A vssd1 vssd1 vccd1 vccd1 _8099_/A sky130_fd_sc_hd__clkbuf_2
X_5897_ _5897_/A _5897_/B vssd1 vssd1 vccd1 vccd1 _5975_/B sky130_fd_sc_hd__xnor2_1
X_4917_ _4917_/A _5066_/B vssd1 vssd1 vccd1 vccd1 _5183_/A sky130_fd_sc_hd__nand2_1
X_8685_ _8704_/CLK _8685_/D vssd1 vssd1 vccd1 vccd1 _8685_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7636_ _7637_/A _7637_/B vssd1 vssd1 vccd1 vccd1 _7638_/A sky130_fd_sc_hd__nor2_1
X_4848_ _4947_/A vssd1 vssd1 vccd1 vccd1 _4851_/A sky130_fd_sc_hd__inv_2
XFILLER_32_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4779_ _4549_/A _5313_/B _4861_/B _4767_/B vssd1 vssd1 vccd1 vccd1 _4779_/X sky130_fd_sc_hd__a22o_1
X_7567_ _8762_/Q _7579_/B vssd1 vssd1 vccd1 vccd1 _7569_/A sky130_fd_sc_hd__xnor2_1
XFILLER_4_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7498_ _7498_/A _7498_/B vssd1 vssd1 vccd1 vccd1 _7499_/B sky130_fd_sc_hd__xnor2_1
X_6518_ _6518_/A vssd1 vssd1 vccd1 vccd1 _8742_/D sky130_fd_sc_hd__clkbuf_1
X_6449_ _8743_/Q _6448_/X _8744_/Q vssd1 vssd1 vccd1 vccd1 _6450_/B sky130_fd_sc_hd__a21o_1
X_8119_ _8119_/A _8038_/B vssd1 vssd1 vccd1 vccd1 _8131_/A sky130_fd_sc_hd__or2b_1
XFILLER_0_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8840__57 vssd1 vssd1 vccd1 vccd1 _8840__57/HI _8949_/A sky130_fd_sc_hd__conb_1
XFILLER_62_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5820_ _5986_/B _5820_/B _5890_/A vssd1 vssd1 vccd1 vccd1 _5890_/B sky130_fd_sc_hd__nand3_1
XFILLER_62_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5751_ _5751_/A vssd1 vssd1 vccd1 vccd1 _6004_/B sky130_fd_sc_hd__clkbuf_2
X_8470_ _8470_/A _8470_/B vssd1 vssd1 vccd1 vccd1 _8471_/B sky130_fd_sc_hd__nor2_1
X_4702_ _4702_/A _4702_/B _4702_/C _4702_/D vssd1 vssd1 vccd1 vccd1 _4771_/B sky130_fd_sc_hd__or4_1
X_5682_ _6147_/A _5682_/B vssd1 vssd1 vccd1 vccd1 _6149_/C sky130_fd_sc_hd__nand2_1
X_7421_ _6910_/C _7285_/B _7420_/Y _7287_/B vssd1 vssd1 vccd1 vccd1 _7487_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_30_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4633_ _4637_/C _4633_/B vssd1 vssd1 vccd1 vccd1 _8635_/D sky130_fd_sc_hd__nor2_1
X_7352_ _7352_/A _7341_/A vssd1 vssd1 vccd1 vccd1 _7352_/X sky130_fd_sc_hd__or2b_1
X_4564_ _4555_/X _4558_/X _4563_/X _5181_/A vssd1 vssd1 vccd1 vccd1 _4566_/B sky130_fd_sc_hd__o31a_1
X_6303_ _6303_/A _6303_/B vssd1 vssd1 vccd1 vccd1 _6304_/B sky130_fd_sc_hd__xnor2_1
X_7283_ _7123_/B _6910_/C _7185_/A _7274_/A vssd1 vssd1 vccd1 vccd1 _7406_/A sky130_fd_sc_hd__a22oi_2
X_6234_ _6234_/A _6234_/B vssd1 vssd1 vccd1 vccd1 _6237_/A sky130_fd_sc_hd__xnor2_1
XFILLER_89_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4495_ _8658_/Q vssd1 vssd1 vccd1 vccd1 _6660_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_103_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6165_ _6166_/A _6165_/B vssd1 vssd1 vccd1 vccd1 _6173_/A sky130_fd_sc_hd__nor2_2
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6096_ _6203_/B _6096_/B vssd1 vssd1 vccd1 vccd1 _6190_/B sky130_fd_sc_hd__nand2_1
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5116_ _5116_/A _5116_/B vssd1 vssd1 vccd1 vccd1 _5116_/X sky130_fd_sc_hd__or2_1
XFILLER_69_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5047_ _5047_/A vssd1 vssd1 vccd1 vccd1 _5255_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_38_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6998_ _6920_/A _7000_/B _6919_/B _6940_/A _6940_/B vssd1 vssd1 vccd1 vccd1 _7165_/A
+ sky130_fd_sc_hd__a32o_1
XFILLER_25_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5949_ _5950_/A _5950_/B vssd1 vssd1 vccd1 vccd1 _6044_/A sky130_fd_sc_hd__nand2_2
XFILLER_25_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8737_ _8742_/CLK _8737_/D vssd1 vssd1 vccd1 vccd1 _8737_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8668_ _8758_/CLK _8668_/D vssd1 vssd1 vccd1 vccd1 _8668_/Q sky130_fd_sc_hd__dfxtp_1
X_8599_ _8599_/A _8612_/B vssd1 vssd1 vccd1 vccd1 _8600_/B sky130_fd_sc_hd__and2_1
X_7619_ _7665_/A _7619_/B _7619_/C _7619_/D vssd1 vssd1 vccd1 vccd1 _7619_/X sky130_fd_sc_hd__or4_1
XFILLER_68_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7970_ _7970_/A _7970_/B vssd1 vssd1 vccd1 vccd1 _7971_/B sky130_fd_sc_hd__nand2_1
XFILLER_66_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6921_ _6802_/A _6885_/A _6886_/B _6814_/A vssd1 vssd1 vccd1 vccd1 _6939_/A sky130_fd_sc_hd__a2bb2o_1
X_6852_ _6757_/A _6757_/B _6757_/C _6851_/Y _6769_/A vssd1 vssd1 vccd1 vccd1 _7011_/A
+ sky130_fd_sc_hd__o311a_2
XFILLER_35_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5803_ _5803_/A _5803_/B vssd1 vssd1 vccd1 vccd1 _5804_/B sky130_fd_sc_hd__or2_1
XFILLER_22_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8522_ _8467_/A _8520_/X _8521_/X vssd1 vssd1 vccd1 vccd1 _8526_/A sky130_fd_sc_hd__a21o_1
X_6783_ _6840_/A _6840_/B vssd1 vssd1 vccd1 vccd1 _6788_/A sky130_fd_sc_hd__xnor2_1
X_5734_ _5993_/A vssd1 vssd1 vccd1 vccd1 _6081_/A sky130_fd_sc_hd__clkinv_2
XFILLER_13_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8453_ _8453_/A _8517_/B vssd1 vssd1 vccd1 vccd1 _8528_/B sky130_fd_sc_hd__xnor2_2
X_5665_ _5764_/A _5796_/B vssd1 vssd1 vccd1 vccd1 _5666_/B sky130_fd_sc_hd__xnor2_1
XFILLER_30_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8384_ _8384_/A _8459_/B _8384_/C vssd1 vssd1 vccd1 vccd1 _8387_/A sky130_fd_sc_hd__nand3_1
X_7404_ _7268_/A _7501_/A _7266_/C _7403_/X vssd1 vssd1 vccd1 vccd1 _7497_/A sky130_fd_sc_hd__a22o_1
X_4616_ _8631_/Q _4616_/B vssd1 vssd1 vccd1 vccd1 _8631_/D sky130_fd_sc_hd__nor2_1
X_5596_ _6378_/D _5645_/C _5595_/Y vssd1 vssd1 vccd1 vccd1 _5597_/B sky130_fd_sc_hd__o21a_1
X_7335_ _7335_/A _7335_/B vssd1 vssd1 vccd1 vccd1 _7356_/B sky130_fd_sc_hd__xor2_1
XFILLER_104_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4547_ _8670_/Q vssd1 vssd1 vccd1 vccd1 _4814_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_4478_ _4480_/A vssd1 vssd1 vccd1 vccd1 _4478_/Y sky130_fd_sc_hd__inv_2
XFILLER_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7266_ _7274_/A _7266_/B _7266_/C vssd1 vssd1 vccd1 vccd1 _7268_/B sky130_fd_sc_hd__nand3_1
X_6217_ _6214_/B _6217_/B vssd1 vssd1 vccd1 vccd1 _6290_/A sky130_fd_sc_hd__and2b_1
X_7197_ _7212_/A _7040_/B _7196_/X vssd1 vssd1 vccd1 vccd1 _7216_/A sky130_fd_sc_hd__o21ai_1
X_6148_ _6149_/C _6227_/A _5527_/A vssd1 vssd1 vccd1 vccd1 _6150_/B sky130_fd_sc_hd__a21o_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_12 _8985_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6079_ _5620_/A _5619_/B _5620_/B _5739_/Y _5979_/A vssd1 vssd1 vccd1 vccd1 _6194_/A
+ sky130_fd_sc_hd__o311a_2
XFILLER_85_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8810__27 vssd1 vssd1 vccd1 vccd1 _8810__27/HI _8905_/A sky130_fd_sc_hd__conb_1
XFILLER_63_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5450_ _5450_/A vssd1 vssd1 vccd1 vccd1 _5450_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4401_ input1/X vssd1 vssd1 vccd1 vccd1 _4426_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5381_ _8694_/Q _5381_/B vssd1 vssd1 vccd1 vccd1 _5387_/C sky130_fd_sc_hd__and2_1
Xclkbuf_3_2_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_5_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7120_ _7120_/A _7120_/B vssd1 vssd1 vccd1 vccd1 _7134_/A sky130_fd_sc_hd__nor2_1
XFILLER_99_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7051_ _7205_/B _7229_/A _7004_/B _7050_/A vssd1 vssd1 vccd1 vccd1 _7052_/B sky130_fd_sc_hd__a2bb2o_1
X_6002_ _6002_/A _5977_/B vssd1 vssd1 vccd1 vccd1 _6007_/A sky130_fd_sc_hd__or2b_1
XFILLER_39_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7953_ _7940_/C _7855_/B _7783_/A _8293_/A vssd1 vssd1 vccd1 vccd1 _7955_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_54_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6904_ _7001_/A _6904_/B vssd1 vssd1 vccd1 vccd1 _6905_/B sky130_fd_sc_hd__xnor2_1
X_7884_ _7888_/A _7888_/B vssd1 vssd1 vccd1 vccd1 _7889_/A sky130_fd_sc_hd__nand2_1
XFILLER_23_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6835_ _6835_/A vssd1 vssd1 vccd1 vccd1 _6910_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_23_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6766_ _6778_/B _6793_/C vssd1 vssd1 vccd1 vccd1 _6767_/C sky130_fd_sc_hd__xnor2_1
X_8505_ _8505_/A _8505_/B vssd1 vssd1 vccd1 vccd1 _8538_/A sky130_fd_sc_hd__xnor2_1
X_5717_ _6068_/A _6378_/D _5717_/C vssd1 vssd1 vccd1 vccd1 _5717_/X sky130_fd_sc_hd__and3_1
X_6697_ _7002_/C vssd1 vssd1 vccd1 vccd1 _7205_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_8436_ _8434_/Y _8401_/B _8435_/Y vssd1 vssd1 vccd1 vccd1 _8472_/A sky130_fd_sc_hd__a21o_1
X_5648_ _5648_/A _8671_/Q vssd1 vssd1 vccd1 vccd1 _5925_/A sky130_fd_sc_hd__nand2_1
X_8367_ _8439_/A _8270_/B _8389_/B _7745_/A vssd1 vssd1 vccd1 vccd1 _8369_/B sky130_fd_sc_hd__a22o_1
X_5579_ _5680_/A _5584_/B vssd1 vssd1 vccd1 vccd1 _5687_/A sky130_fd_sc_hd__nand2_2
X_8298_ _8299_/A _8299_/B vssd1 vssd1 vccd1 vccd1 _8345_/A sky130_fd_sc_hd__nor2_1
X_8876__93 vssd1 vssd1 vccd1 vccd1 _8876__93/HI _8985_/A sky130_fd_sc_hd__conb_1
X_7318_ _7318_/A _7318_/B _7318_/C vssd1 vssd1 vccd1 vccd1 _7319_/B sky130_fd_sc_hd__and3_1
X_7249_ _7068_/A _7248_/B _7248_/A vssd1 vssd1 vccd1 vccd1 _7249_/X sky130_fd_sc_hd__o21ba_1
XFILLER_104_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4950_ _5251_/B vssd1 vssd1 vccd1 vccd1 _4950_/X sky130_fd_sc_hd__clkbuf_2
X_4881_ _4850_/C _4927_/B _4874_/B vssd1 vssd1 vccd1 vccd1 _4882_/B sky130_fd_sc_hd__a21oi_1
XFILLER_32_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6620_ _6621_/B _8748_/Q vssd1 vssd1 vccd1 vccd1 _6645_/A sky130_fd_sc_hd__nand2b_2
X_6551_ _8751_/Q vssd1 vssd1 vccd1 vccd1 _6583_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5502_ _5500_/X _5505_/A vssd1 vssd1 vccd1 vccd1 _5547_/B sky130_fd_sc_hd__and2b_1
X_6482_ _6482_/A _6486_/C vssd1 vssd1 vccd1 vccd1 _6485_/A sky130_fd_sc_hd__and2_1
X_8221_ _8221_/A _8221_/B vssd1 vssd1 vccd1 vccd1 _8222_/B sky130_fd_sc_hd__nand2_1
X_5433_ _8710_/Q vssd1 vssd1 vccd1 vccd1 _5463_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_8152_ _8080_/A _8080_/B _8151_/Y vssd1 vssd1 vccd1 vccd1 _8180_/A sky130_fd_sc_hd__o21a_2
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5364_ _6532_/B _5365_/C _5363_/Y vssd1 vssd1 vccd1 vccd1 _8688_/D sky130_fd_sc_hd__a21oi_1
X_7103_ _7104_/A _7104_/B vssd1 vssd1 vccd1 vccd1 _7108_/A sky130_fd_sc_hd__or2b_1
X_8083_ _8083_/A _8013_/B vssd1 vssd1 vccd1 vccd1 _8083_/X sky130_fd_sc_hd__or2b_1
X_5295_ _5271_/X _5294_/X _4974_/X vssd1 vssd1 vccd1 vccd1 _5296_/D sky130_fd_sc_hd__a21oi_1
XFILLER_87_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7034_ _7034_/A _7034_/B vssd1 vssd1 vccd1 vccd1 _7035_/A sky130_fd_sc_hd__nor2_1
XFILLER_19_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8985_ _8985_/A _4482_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[34] sky130_fd_sc_hd__ebufn_8
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7936_ _7981_/A _7981_/B _7981_/C vssd1 vssd1 vccd1 vccd1 _7964_/A sky130_fd_sc_hd__nand3_1
X_7867_ _7867_/A _7893_/A _7867_/C vssd1 vssd1 vccd1 vccd1 _7976_/A sky130_fd_sc_hd__or3_1
X_6818_ _6818_/A _6818_/B vssd1 vssd1 vccd1 vccd1 _6820_/B sky130_fd_sc_hd__or2_1
XFILLER_23_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7798_ _7924_/A _7826_/A vssd1 vssd1 vccd1 vccd1 _7818_/A sky130_fd_sc_hd__nand2_1
XFILLER_51_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6749_ _6793_/A _7080_/C vssd1 vssd1 vccd1 vccd1 _7119_/A sky130_fd_sc_hd__nor2_1
X_8419_ _8418_/Y _8351_/B _8349_/X vssd1 vssd1 vccd1 vccd1 _8421_/A sky130_fd_sc_hd__a21boi_1
XFILLER_104_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5080_ _5172_/C _5261_/D vssd1 vssd1 vccd1 vccd1 _5149_/D sky130_fd_sc_hd__or2_1
XFILLER_96_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5982_ _6183_/B _5893_/X _5892_/Y _6193_/A vssd1 vssd1 vccd1 vccd1 _6088_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_64_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8770_ _8784_/CLK _8770_/D vssd1 vssd1 vccd1 vccd1 _8770_/Q sky130_fd_sc_hd__dfxtp_1
X_7721_ _6655_/B _8783_/Q vssd1 vssd1 vccd1 vccd1 _7722_/B sky130_fd_sc_hd__and2b_1
XFILLER_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4933_ _5062_/A _4942_/A vssd1 vssd1 vccd1 vccd1 _5201_/A sky130_fd_sc_hd__or2_4
X_7652_ _7640_/B _7652_/B _7652_/C vssd1 vssd1 vccd1 vccd1 _7652_/X sky130_fd_sc_hd__and3b_1
X_4864_ _5053_/B _5266_/B vssd1 vssd1 vccd1 vccd1 _5123_/A sky130_fd_sc_hd__nand2_1
X_7583_ _7583_/A _7583_/B vssd1 vssd1 vccd1 vccd1 _7583_/Y sky130_fd_sc_hd__nand2_1
XFILLER_32_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4795_ _5501_/B _4796_/B vssd1 vssd1 vccd1 vccd1 _4804_/C sky130_fd_sc_hd__nor2_1
X_6603_ _6593_/A _6590_/C _6597_/D _6602_/X vssd1 vssd1 vccd1 vccd1 _6604_/C sky130_fd_sc_hd__o31a_1
X_6534_ _6534_/A _6534_/B _6534_/C vssd1 vssd1 vccd1 vccd1 _6535_/D sky130_fd_sc_hd__or3_1
XFILLER_21_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6465_ _6517_/B vssd1 vssd1 vccd1 vccd1 _6465_/X sky130_fd_sc_hd__clkbuf_2
X_8204_ _8204_/A _8204_/B vssd1 vssd1 vccd1 vccd1 _8205_/B sky130_fd_sc_hd__nor2_1
X_5416_ _8719_/Q vssd1 vssd1 vccd1 vccd1 _6405_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6396_ _8574_/A _8716_/Q vssd1 vssd1 vccd1 vccd1 _6396_/Y sky130_fd_sc_hd__nor2_1
X_8846__63 vssd1 vssd1 vccd1 vccd1 _8846__63/HI _8955_/A sky130_fd_sc_hd__conb_1
XFILLER_99_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8135_ _8135_/A _8135_/B vssd1 vssd1 vccd1 vccd1 _8311_/B sky130_fd_sc_hd__xor2_2
X_5347_ _5355_/A vssd1 vssd1 vccd1 vccd1 _6567_/A sky130_fd_sc_hd__buf_2
XFILLER_87_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8066_ _7996_/A _8155_/B _8155_/C _8258_/A vssd1 vssd1 vccd1 vccd1 _8066_/X sky130_fd_sc_hd__a31o_1
X_5278_ _5278_/A _5278_/B _5278_/C vssd1 vssd1 vccd1 vccd1 _5278_/X sky130_fd_sc_hd__or3_1
XFILLER_75_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7017_ _6914_/A _7017_/B vssd1 vssd1 vccd1 vccd1 _7017_/X sky130_fd_sc_hd__and2b_1
XFILLER_68_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8968_ _8968_/A _4461_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[17] sky130_fd_sc_hd__ebufn_8
XFILLER_43_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7919_ _7919_/A _7919_/B _7919_/C vssd1 vssd1 vccd1 vccd1 _7921_/B sky130_fd_sc_hd__nand3_1
XFILLER_15_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8899_ _8899_/A _4380_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[18] sky130_fd_sc_hd__ebufn_8
XFILLER_70_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4580_ _8674_/Q _4584_/B vssd1 vssd1 vccd1 vccd1 _4581_/A sky130_fd_sc_hd__and2_2
XFILLER_52_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6250_ _6250_/A _6251_/B _6311_/C vssd1 vssd1 vccd1 vccd1 _6337_/A sky130_fd_sc_hd__and3_1
X_6181_ _6181_/A _6181_/B vssd1 vssd1 vccd1 vccd1 _6181_/Y sky130_fd_sc_hd__nand2_1
X_5201_ _5201_/A _5201_/B _5228_/B vssd1 vssd1 vccd1 vccd1 _5227_/B sky130_fd_sc_hd__or3_1
X_5132_ _4977_/A _5131_/X _5296_/A vssd1 vssd1 vccd1 vccd1 _5132_/X sky130_fd_sc_hd__o21ba_1
XFILLER_96_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5063_ _5250_/D _5163_/C _5211_/A _5128_/A vssd1 vssd1 vccd1 vccd1 _5071_/C sky130_fd_sc_hd__or4_1
XFILLER_37_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5965_ _5965_/A _6370_/A _5965_/C vssd1 vssd1 vccd1 vccd1 _5965_/Y sky130_fd_sc_hd__nor3_1
XFILLER_80_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8753_ _8753_/CLK _8753_/D vssd1 vssd1 vccd1 vccd1 _8753_/Q sky130_fd_sc_hd__dfxtp_1
X_7704_ _8354_/A vssd1 vssd1 vccd1 vccd1 _8293_/A sky130_fd_sc_hd__clkbuf_2
X_5896_ _5977_/A _5977_/B vssd1 vssd1 vccd1 vccd1 _5897_/B sky130_fd_sc_hd__xor2_1
XFILLER_21_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4916_ _5009_/C _4916_/B vssd1 vssd1 vccd1 vccd1 _5066_/B sky130_fd_sc_hd__nand2_2
X_8684_ _8704_/CLK _8684_/D vssd1 vssd1 vccd1 vccd1 _8684_/Q sky130_fd_sc_hd__dfxtp_1
X_7635_ _7630_/A _7627_/X _7634_/X _5335_/X vssd1 vssd1 vccd1 vccd1 _8769_/D sky130_fd_sc_hd__o211a_1
X_4847_ _4938_/A vssd1 vssd1 vccd1 vccd1 _5159_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_32_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4778_ _4778_/A _4850_/A vssd1 vssd1 vccd1 vccd1 _4861_/B sky130_fd_sc_hd__nand2_1
X_7566_ _7562_/A _6567_/X _6569_/A _7565_/X vssd1 vssd1 vccd1 vccd1 _8761_/D sky130_fd_sc_hd__a22o_1
X_7497_ _7497_/A _7497_/B vssd1 vssd1 vccd1 vccd1 _7498_/B sky130_fd_sc_hd__xnor2_1
X_6517_ _6519_/B _6517_/B _6517_/C vssd1 vssd1 vccd1 vccd1 _6518_/A sky130_fd_sc_hd__and3b_1
X_6448_ _8740_/Q _6515_/B _6456_/B _6447_/X _8742_/Q vssd1 vssd1 vccd1 vccd1 _6448_/X
+ sky130_fd_sc_hd__a221o_1
X_6379_ _6381_/A _6377_/X _6378_/X vssd1 vssd1 vccd1 vccd1 _6388_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8118_ _8145_/B _8118_/B vssd1 vssd1 vccd1 vccd1 _8133_/A sky130_fd_sc_hd__xnor2_1
XFILLER_87_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8049_ _7972_/A _7974_/A _8057_/B _8048_/X vssd1 vssd1 vccd1 vccd1 _8055_/A sky130_fd_sc_hd__o211a_1
XFILLER_87_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5750_ _6004_/A _5824_/B _5750_/C vssd1 vssd1 vccd1 vccd1 _5754_/B sky130_fd_sc_hd__and3_1
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5681_ _5681_/A _6378_/B vssd1 vssd1 vccd1 vccd1 _5697_/A sky130_fd_sc_hd__nand2_1
X_4701_ _4701_/A vssd1 vssd1 vccd1 vccd1 _4702_/D sky130_fd_sc_hd__clkbuf_2
X_7420_ _7420_/A vssd1 vssd1 vccd1 vccd1 _7420_/Y sky130_fd_sc_hd__clkinv_2
X_4632_ _8635_/Q _4630_/A _4628_/X vssd1 vssd1 vccd1 vccd1 _4633_/B sky130_fd_sc_hd__o21ai_1
X_7351_ _7344_/A _7344_/B _7350_/Y vssd1 vssd1 vccd1 vccd1 _7433_/A sky130_fd_sc_hd__a21o_1
X_4563_ _5263_/A vssd1 vssd1 vccd1 vccd1 _4563_/X sky130_fd_sc_hd__clkbuf_2
X_6302_ _6302_/A _6302_/B vssd1 vssd1 vccd1 vccd1 _6303_/B sky130_fd_sc_hd__xnor2_1
X_7282_ _7282_/A _7282_/B vssd1 vssd1 vccd1 vccd1 _7284_/A sky130_fd_sc_hd__xor2_1
X_4494_ _6613_/B vssd1 vssd1 vccd1 vccd1 _5181_/A sky130_fd_sc_hd__clkbuf_2
X_6233_ _6233_/A _6307_/B vssd1 vssd1 vccd1 vccd1 _6234_/B sky130_fd_sc_hd__xnor2_1
XFILLER_6_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8816__33 vssd1 vssd1 vccd1 vccd1 _8816__33/HI _8911_/A sky130_fd_sc_hd__conb_1
X_6164_ _6104_/A _6104_/B _6163_/X vssd1 vssd1 vccd1 vccd1 _6212_/A sky130_fd_sc_hd__a21oi_1
XFILLER_69_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6095_ _6095_/A _6277_/B vssd1 vssd1 vccd1 vccd1 _6096_/B sky130_fd_sc_hd__nand2_1
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5115_ _5163_/C _5263_/C _5206_/B _5188_/D vssd1 vssd1 vccd1 vccd1 _5116_/B sky130_fd_sc_hd__or4_1
XFILLER_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5046_ _4733_/B _5281_/A _5018_/X _5045_/X _4819_/A vssd1 vssd1 vccd1 vccd1 _5073_/A
+ sky130_fd_sc_hd__o311a_1
XFILLER_72_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6997_ _6954_/A _6954_/B _6996_/X vssd1 vssd1 vccd1 vccd1 _7062_/A sky130_fd_sc_hd__a21o_1
X_5948_ _6121_/A _5948_/B vssd1 vssd1 vccd1 vccd1 _5950_/B sky130_fd_sc_hd__nor2_1
XFILLER_53_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8736_ _8742_/CLK _8736_/D vssd1 vssd1 vccd1 vccd1 _8736_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5879_ _5879_/A _5883_/A _5879_/C vssd1 vssd1 vccd1 vccd1 _5881_/B sky130_fd_sc_hd__or3_1
X_8667_ _8771_/CLK _8667_/D vssd1 vssd1 vccd1 vccd1 _8667_/Q sky130_fd_sc_hd__dfxtp_1
X_8598_ _8599_/A _8612_/B vssd1 vssd1 vccd1 vccd1 _8600_/A sky130_fd_sc_hd__nor2_1
X_7618_ _7637_/A _7630_/A _7649_/A vssd1 vssd1 vccd1 vccd1 _7619_/D sky130_fd_sc_hd__o21a_1
XFILLER_21_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7549_ _7551_/B _7548_/Y _7552_/A _7552_/B vssd1 vssd1 vccd1 vccd1 _7549_/X sky130_fd_sc_hd__a211o_1
XFILLER_68_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_4_0_wb_clk_i clkbuf_4_5_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _8730_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_16_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6920_ _6920_/A _6920_/B vssd1 vssd1 vccd1 vccd1 _6940_/A sky130_fd_sc_hd__xor2_1
XFILLER_47_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6851_ _6851_/A _8671_/Q vssd1 vssd1 vccd1 vccd1 _6851_/Y sky130_fd_sc_hd__nand2_1
X_5802_ _5801_/A _5801_/B _5801_/C vssd1 vssd1 vccd1 vccd1 _5803_/B sky130_fd_sc_hd__o21a_1
X_8521_ _8521_/A _8521_/B vssd1 vssd1 vccd1 vccd1 _8521_/X sky130_fd_sc_hd__and2_1
XFILLER_22_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6782_ _7118_/A _7020_/A _6782_/C vssd1 vssd1 vccd1 vccd1 _6840_/B sky130_fd_sc_hd__and3_1
X_5733_ _5991_/A _6192_/A vssd1 vssd1 vccd1 vccd1 _5743_/A sky130_fd_sc_hd__nor2_1
X_8452_ _8452_/A _8516_/B vssd1 vssd1 vccd1 vccd1 _8517_/B sky130_fd_sc_hd__xnor2_1
X_5664_ _5766_/C _5664_/B vssd1 vssd1 vccd1 vccd1 _5796_/B sky130_fd_sc_hd__xor2_1
XFILLER_30_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8383_ _8380_/X _8459_/A _8263_/B vssd1 vssd1 vccd1 vccd1 _8384_/C sky130_fd_sc_hd__a21o_1
X_5595_ _5984_/C _5701_/B _6262_/B vssd1 vssd1 vccd1 vccd1 _5595_/Y sky130_fd_sc_hd__nand3_2
X_4615_ _4615_/A _5443_/B vssd1 vssd1 vccd1 vccd1 _4616_/B sky130_fd_sc_hd__nand2_2
X_7403_ _7411_/A _7411_/B _7268_/B vssd1 vssd1 vccd1 vccd1 _7403_/X sky130_fd_sc_hd__o21a_1
X_7334_ _7334_/A _7370_/C vssd1 vssd1 vccd1 vccd1 _7335_/B sky130_fd_sc_hd__xnor2_1
X_4546_ _6758_/B _4568_/B _4543_/Y _7943_/B vssd1 vssd1 vccd1 vccd1 _4574_/A sky130_fd_sc_hd__o31a_1
X_4477_ _4480_/A vssd1 vssd1 vccd1 vccd1 _4477_/Y sky130_fd_sc_hd__inv_2
X_7265_ _7279_/A _7279_/B _7265_/C vssd1 vssd1 vccd1 vccd1 _7266_/C sky130_fd_sc_hd__or3_1
X_6216_ _6294_/A _6294_/B vssd1 vssd1 vccd1 vccd1 _6292_/A sky130_fd_sc_hd__nand2_1
X_7196_ _7196_/A _7039_/A vssd1 vssd1 vccd1 vccd1 _7196_/X sky130_fd_sc_hd__or2b_1
X_6147_ _6147_/A _6169_/B vssd1 vssd1 vccd1 vccd1 _6227_/A sky130_fd_sc_hd__or2_1
XFILLER_57_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_13 _8985_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6078_ _6000_/A _6075_/B _5999_/B _6077_/Y vssd1 vssd1 vccd1 vccd1 _6101_/A sky130_fd_sc_hd__o31ai_4
XFILLER_57_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5029_ _5042_/D vssd1 vssd1 vccd1 vccd1 _5128_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_26_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8719_ _8720_/CLK _8719_/D vssd1 vssd1 vccd1 vccd1 _8719_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_9_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4400_ _4400_/A vssd1 vssd1 vccd1 vccd1 _4400_/Y sky130_fd_sc_hd__inv_2
X_5380_ _5380_/A vssd1 vssd1 vccd1 vccd1 _8693_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7050_ _7050_/A _7392_/B vssd1 vssd1 vccd1 vccd1 _7227_/A sky130_fd_sc_hd__nor2_1
XFILLER_86_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6001_ _6001_/A _6066_/B vssd1 vssd1 vccd1 vccd1 _6009_/A sky130_fd_sc_hd__xnor2_2
XFILLER_67_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7952_ _8036_/A _8036_/B vssd1 vssd1 vccd1 vccd1 _7958_/A sky130_fd_sc_hd__xnor2_1
XFILLER_54_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6903_ _7282_/A _7416_/B _7022_/A vssd1 vssd1 vccd1 vccd1 _6904_/B sky130_fd_sc_hd__a21oi_2
X_7883_ _8567_/A _8567_/B _8571_/B vssd1 vssd1 vccd1 vccd1 _7888_/B sky130_fd_sc_hd__and3_1
XFILLER_62_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6834_ _7198_/B _6834_/B vssd1 vssd1 vccd1 vccd1 _6848_/A sky130_fd_sc_hd__xnor2_1
XFILLER_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6765_ _6765_/A _6910_/B vssd1 vssd1 vccd1 vccd1 _6793_/C sky130_fd_sc_hd__nand2_1
X_8504_ _8471_/A _8470_/B _8470_/A vssd1 vssd1 vccd1 vccd1 _8505_/B sky130_fd_sc_hd__o21bai_1
X_5716_ _5643_/A _5716_/B vssd1 vssd1 vccd1 vccd1 _5810_/A sky130_fd_sc_hd__and2b_1
X_8435_ _8435_/A _8435_/B vssd1 vssd1 vccd1 vccd1 _8435_/Y sky130_fd_sc_hd__nor2_1
X_6696_ _6696_/A _6696_/B vssd1 vssd1 vccd1 vccd1 _7002_/C sky130_fd_sc_hd__xor2_2
X_5647_ _5512_/B _6142_/B _5531_/D _5556_/A vssd1 vssd1 vccd1 vccd1 _5764_/A sky130_fd_sc_hd__o31a_1
XFILLER_40_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8366_ _8268_/A _8268_/C _8268_/B vssd1 vssd1 vccd1 vccd1 _8438_/B sky130_fd_sc_hd__a21bo_1
X_5578_ _6402_/S _7739_/B vssd1 vssd1 vccd1 vccd1 _5584_/B sky130_fd_sc_hd__nand2_1
XFILLER_104_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8297_ _8124_/B _8216_/B _8214_/Y vssd1 vssd1 vccd1 vccd1 _8299_/B sky130_fd_sc_hd__a21o_1
X_7317_ _7318_/A _7318_/B _7318_/C vssd1 vssd1 vccd1 vccd1 _7319_/A sky130_fd_sc_hd__a21oi_1
XFILLER_2_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4529_ _7775_/B vssd1 vssd1 vccd1 vccd1 _6758_/B sky130_fd_sc_hd__buf_2
X_7248_ _7248_/A _7248_/B vssd1 vssd1 vccd1 vccd1 _7533_/A sky130_fd_sc_hd__nor2_1
XFILLER_77_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7179_ _7179_/A _7179_/B vssd1 vssd1 vccd1 vccd1 _7180_/B sky130_fd_sc_hd__or2_1
XFILLER_100_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4880_ _4934_/A _4894_/B _4915_/B _4879_/X vssd1 vssd1 vccd1 vccd1 _5261_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6550_ _8749_/Q vssd1 vssd1 vccd1 vccd1 _6570_/A sky130_fd_sc_hd__clkbuf_2
X_5501_ _8709_/Q _5501_/B vssd1 vssd1 vccd1 vccd1 _5505_/A sky130_fd_sc_hd__nand2_2
XFILLER_9_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6481_ _6481_/A vssd1 vssd1 vccd1 vccd1 _8730_/D sky130_fd_sc_hd__clkbuf_1
X_8220_ _8220_/A _8220_/B vssd1 vssd1 vccd1 vccd1 _8221_/B sky130_fd_sc_hd__or2_1
X_5432_ _8708_/Q vssd1 vssd1 vccd1 vccd1 _5452_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_99_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8151_ _8151_/A _8151_/B vssd1 vssd1 vccd1 vccd1 _8151_/Y sky130_fd_sc_hd__nand2_1
X_5363_ _6532_/B _5365_/C _5409_/A vssd1 vssd1 vccd1 vccd1 _5363_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_99_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7102_ _6782_/C _7101_/Y _6961_/B vssd1 vssd1 vccd1 vccd1 _7104_/B sky130_fd_sc_hd__o21a_1
XFILLER_101_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8082_ _8082_/A _8082_/B vssd1 vssd1 vccd1 vccd1 _8082_/Y sky130_fd_sc_hd__nand2_1
X_5294_ _4702_/C _5269_/A _5279_/X _5293_/X _5170_/A vssd1 vssd1 vccd1 vccd1 _5294_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_101_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7033_ _7019_/A _6912_/B _6910_/X vssd1 vssd1 vccd1 vccd1 _7037_/A sky130_fd_sc_hd__a21oi_2
XFILLER_19_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8984_ _8984_/A _4480_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[33] sky130_fd_sc_hd__ebufn_8
XFILLER_82_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7935_ _7934_/A _7934_/B _7934_/C _7934_/D vssd1 vssd1 vccd1 vccd1 _7981_/C sky130_fd_sc_hd__a22o_1
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7866_ _7866_/A _7866_/B vssd1 vssd1 vccd1 vccd1 _7867_/C sky130_fd_sc_hd__and2_1
XFILLER_23_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6817_ _6816_/A _6949_/A _6729_/A _6729_/B _6726_/Y vssd1 vssd1 vccd1 vccd1 _6818_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_23_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7797_ _7912_/A _7912_/B vssd1 vssd1 vccd1 vccd1 _7826_/A sky130_fd_sc_hd__xor2_2
XFILLER_23_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6748_ _6784_/B vssd1 vssd1 vccd1 vccd1 _7080_/C sky130_fd_sc_hd__clkbuf_2
X_6679_ _6679_/A _6679_/B vssd1 vssd1 vccd1 vccd1 _6688_/A sky130_fd_sc_hd__xor2_2
X_8418_ _8418_/A vssd1 vssd1 vccd1 vccd1 _8418_/Y sky130_fd_sc_hd__inv_2
X_8349_ _8349_/A _8498_/S vssd1 vssd1 vccd1 vccd1 _8349_/X sky130_fd_sc_hd__or2_1
XFILLER_104_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5981_ _6068_/B _5981_/B vssd1 vssd1 vccd1 vccd1 _5988_/A sky130_fd_sc_hd__xnor2_2
XFILLER_52_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7720_ _8783_/Q _8659_/Q vssd1 vssd1 vccd1 vccd1 _7722_/A sky130_fd_sc_hd__and2b_2
XFILLER_52_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4932_ _5077_/B _5251_/A vssd1 vssd1 vccd1 vccd1 _4942_/A sky130_fd_sc_hd__or2_1
X_7651_ _7665_/A _7651_/B vssd1 vssd1 vccd1 vccd1 _7654_/B sky130_fd_sc_hd__nand2_1
XFILLER_60_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4863_ _5083_/A _5082_/B vssd1 vssd1 vccd1 vccd1 _5266_/B sky130_fd_sc_hd__or2_2
X_6602_ _6602_/A _6602_/B vssd1 vssd1 vccd1 vccd1 _6602_/X sky130_fd_sc_hd__or2_1
X_4794_ _6627_/B vssd1 vssd1 vccd1 vccd1 _5501_/B sky130_fd_sc_hd__clkinv_2
XFILLER_20_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7582_ _7578_/Y _7586_/S _7579_/Y _7585_/B _7583_/B vssd1 vssd1 vccd1 vccd1 _7582_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_20_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6533_ _8697_/Q _8696_/Q _8704_/Q vssd1 vssd1 vccd1 vccd1 _6534_/C sky130_fd_sc_hd__or3_1
XFILLER_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6464_ _6563_/B _7622_/A vssd1 vssd1 vccd1 vccd1 _6517_/B sky130_fd_sc_hd__and2_1
X_8203_ _8204_/A _8204_/B vssd1 vssd1 vccd1 vccd1 _8302_/B sky130_fd_sc_hd__and2_1
X_5415_ _8720_/Q vssd1 vssd1 vccd1 vccd1 _6409_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6395_ _6398_/B _6394_/Y _6390_/A _6390_/B vssd1 vssd1 vccd1 vccd1 _6395_/X sky130_fd_sc_hd__a211o_1
XFILLER_99_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8134_ _8143_/B _8134_/B vssd1 vssd1 vccd1 vccd1 _8135_/B sky130_fd_sc_hd__xnor2_2
X_5346_ _6563_/B _6562_/A vssd1 vssd1 vccd1 vccd1 _5355_/A sky130_fd_sc_hd__and2_1
XFILLER_87_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8065_ _7813_/A _7807_/B _7813_/C _8381_/A _7754_/A vssd1 vssd1 vccd1 vccd1 _8258_/A
+ sky130_fd_sc_hd__a311oi_4
X_5277_ _5288_/B _5277_/B _5277_/C _5277_/D vssd1 vssd1 vccd1 vccd1 _5278_/C sky130_fd_sc_hd__or4_1
X_8861__78 vssd1 vssd1 vccd1 vccd1 _8861__78/HI _8970_/A sky130_fd_sc_hd__conb_1
XFILLER_87_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7016_ _7169_/A _7016_/B vssd1 vssd1 vccd1 vccd1 _7024_/A sky130_fd_sc_hd__xor2_1
XFILLER_101_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8967_ _8967_/A _4460_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[16] sky130_fd_sc_hd__ebufn_8
X_7918_ _7918_/A _7918_/B vssd1 vssd1 vccd1 vccd1 _7919_/C sky130_fd_sc_hd__xor2_1
X_8898_ _8898_/A _4379_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[17] sky130_fd_sc_hd__ebufn_8
X_7849_ _7859_/A _7940_/C vssd1 vssd1 vccd1 vccd1 _7850_/B sky130_fd_sc_hd__xnor2_1
XFILLER_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6180_ _6183_/A _6180_/B vssd1 vssd1 vccd1 vccd1 _6248_/A sky130_fd_sc_hd__or2_1
X_5200_ _5255_/A _5228_/A _5128_/A _5119_/B _5199_/Y vssd1 vssd1 vccd1 vccd1 _5200_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5131_ _4974_/X _5224_/C _5073_/X _5130_/X vssd1 vssd1 vccd1 vccd1 _5131_/X sky130_fd_sc_hd__o31a_1
X_5062_ _5062_/A vssd1 vssd1 vccd1 vccd1 _5163_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_96_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8752_ _8765_/CLK _8752_/D vssd1 vssd1 vccd1 vccd1 _8752_/Q sky130_fd_sc_hd__dfxtp_1
X_5964_ _6370_/A _6370_/B _6369_/B _6369_/A _6369_/C vssd1 vssd1 vccd1 vccd1 _6367_/B
+ sky130_fd_sc_hd__o2111ai_4
X_7703_ _8190_/A vssd1 vssd1 vccd1 vccd1 _8354_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_80_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5895_ _6183_/B _5895_/B vssd1 vssd1 vccd1 vccd1 _5977_/B sky130_fd_sc_hd__xnor2_2
X_8683_ _8776_/CLK _8683_/D vssd1 vssd1 vccd1 vccd1 _8683_/Q sky130_fd_sc_hd__dfxtp_1
X_4915_ _5009_/C _4915_/B vssd1 vssd1 vccd1 vccd1 _4917_/A sky130_fd_sc_hd__nand2_1
XFILLER_40_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7634_ _8603_/A _7634_/B vssd1 vssd1 vccd1 vccd1 _7634_/X sky130_fd_sc_hd__or2_1
XFILLER_20_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4846_ _5155_/C _5078_/B vssd1 vssd1 vccd1 vccd1 _4938_/A sky130_fd_sc_hd__or2_1
X_7565_ _7565_/A _7565_/B vssd1 vssd1 vccd1 vccd1 _7565_/X sky130_fd_sc_hd__xor2_1
X_4777_ _4897_/B _4765_/X _5313_/B _4877_/C _7606_/A vssd1 vssd1 vccd1 vccd1 _8663_/D
+ sky130_fd_sc_hd__o221a_1
X_6516_ _8740_/Q _6515_/B _6510_/B _8742_/Q vssd1 vssd1 vccd1 vccd1 _6517_/C sky130_fd_sc_hd__a31o_1
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7496_ _7379_/B _6813_/B _7489_/B _6707_/A vssd1 vssd1 vccd1 vccd1 _7497_/B sky130_fd_sc_hd__a22o_1
X_6447_ _8737_/Q _6445_/X _6506_/B vssd1 vssd1 vccd1 vccd1 _6447_/X sky130_fd_sc_hd__a21o_1
X_6378_ _6378_/A _6378_/B _6378_/C _6378_/D vssd1 vssd1 vccd1 vccd1 _6378_/X sky130_fd_sc_hd__and4_1
XFILLER_102_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8117_ _8117_/A _8117_/B vssd1 vssd1 vccd1 vccd1 _8118_/B sky130_fd_sc_hd__xnor2_1
X_5329_ _8755_/Q _5320_/X _5328_/X _5324_/X vssd1 vssd1 vccd1 vccd1 _8680_/D sky130_fd_sc_hd__o211a_1
XFILLER_87_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8048_ _8057_/A _8047_/B _8047_/C vssd1 vssd1 vccd1 vccd1 _8048_/X sky130_fd_sc_hd__a21o_1
XFILLER_102_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8787__4 vssd1 vssd1 vccd1 vccd1 _8787__4/HI _8882_/A sky130_fd_sc_hd__conb_1
XFILLER_98_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5680_ _5680_/A _5680_/B vssd1 vssd1 vccd1 vccd1 _5891_/A sky130_fd_sc_hd__xnor2_2
X_4700_ _5210_/A _5047_/A vssd1 vssd1 vccd1 vccd1 _4701_/A sky130_fd_sc_hd__nand2_1
XFILLER_8_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4631_ _8634_/Q _8635_/Q _4631_/C vssd1 vssd1 vccd1 vccd1 _4637_/C sky130_fd_sc_hd__and3_1
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7350_ _7350_/A _7350_/B vssd1 vssd1 vccd1 vccd1 _7350_/Y sky130_fd_sc_hd__nor2_1
X_4562_ _5138_/A _5066_/A vssd1 vssd1 vccd1 vccd1 _5263_/A sky130_fd_sc_hd__or2_2
X_6301_ _6286_/A _6286_/B _6300_/Y vssd1 vssd1 vccd1 vccd1 _6303_/A sky130_fd_sc_hd__a21bo_1
XFILLER_6_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7281_ _7281_/A _7281_/B vssd1 vssd1 vccd1 vccd1 _7282_/B sky130_fd_sc_hd__xor2_1
X_4493_ _7729_/B vssd1 vssd1 vccd1 vccd1 _6613_/B sky130_fd_sc_hd__buf_2
X_6232_ _6232_/A _6232_/B vssd1 vssd1 vccd1 vccd1 _6307_/B sky130_fd_sc_hd__xor2_1
XFILLER_97_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6163_ _6103_/A _6163_/B vssd1 vssd1 vccd1 vccd1 _6163_/X sky130_fd_sc_hd__and2b_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6094_ _6095_/A _6277_/B vssd1 vssd1 vccd1 vccd1 _6203_/B sky130_fd_sc_hd__or2_1
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5114_ _5172_/A _5288_/C _5119_/B vssd1 vssd1 vccd1 vccd1 _5116_/A sky130_fd_sc_hd__or3_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8831__48 vssd1 vssd1 vccd1 vccd1 _8831__48/HI _8940_/A sky130_fd_sc_hd__conb_1
X_5045_ _5192_/A _5031_/X _5038_/X _5044_/X _4720_/A vssd1 vssd1 vccd1 vccd1 _5045_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_38_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6996_ _6941_/A _6996_/B vssd1 vssd1 vccd1 vccd1 _6996_/X sky130_fd_sc_hd__and2b_1
X_5947_ _5946_/A _5946_/B _5946_/C vssd1 vssd1 vccd1 vccd1 _5948_/B sky130_fd_sc_hd__a21oi_1
XFILLER_80_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8735_ _8742_/CLK _8735_/D vssd1 vssd1 vccd1 vccd1 _8735_/Q sky130_fd_sc_hd__dfxtp_1
X_8666_ _8783_/CLK _8666_/D vssd1 vssd1 vccd1 vccd1 _8666_/Q sky130_fd_sc_hd__dfxtp_4
X_5878_ _5885_/B _5876_/X _5801_/A _5803_/A vssd1 vssd1 vccd1 vccd1 _5879_/C sky130_fd_sc_hd__a211oi_1
X_7617_ _8772_/Q vssd1 vssd1 vccd1 vccd1 _7665_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_8597_ _8593_/A _7627_/X _8596_/X _7642_/X vssd1 vssd1 vccd1 vccd1 _8780_/D sky130_fd_sc_hd__o211a_1
X_4829_ _4927_/A _4927_/B _5298_/C vssd1 vssd1 vccd1 vccd1 _4926_/B sky130_fd_sc_hd__nand3_2
X_7548_ _7548_/A _7548_/B vssd1 vssd1 vccd1 vccd1 _7548_/Y sky130_fd_sc_hd__nand2_1
X_7479_ _7479_/A _7479_/B vssd1 vssd1 vccd1 vccd1 _7480_/B sky130_fd_sc_hd__xnor2_1
XFILLER_68_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6850_ _7301_/A vssd1 vssd1 vccd1 vccd1 _7378_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_35_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5801_ _5801_/A _5801_/B _5801_/C vssd1 vssd1 vccd1 vccd1 _5803_/A sky130_fd_sc_hd__nor3_1
XFILLER_22_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6781_ _6793_/A _7020_/B vssd1 vssd1 vccd1 vccd1 _6782_/C sky130_fd_sc_hd__nor2_1
X_8520_ _8521_/A _8521_/B vssd1 vssd1 vccd1 vccd1 _8520_/X sky130_fd_sc_hd__or2_1
X_5732_ _5732_/A _5732_/B vssd1 vssd1 vccd1 vccd1 _6192_/A sky130_fd_sc_hd__xnor2_2
X_8451_ _8449_/X _8450_/X _8514_/B vssd1 vssd1 vccd1 vccd1 _8516_/B sky130_fd_sc_hd__a21oi_1
X_5663_ _5512_/B _5531_/D _5662_/X vssd1 vssd1 vccd1 vccd1 _5664_/B sky130_fd_sc_hd__o21a_1
X_8382_ _8382_/A _8382_/B vssd1 vssd1 vccd1 vccd1 _8459_/A sky130_fd_sc_hd__nand2_1
X_5594_ _5594_/A vssd1 vssd1 vccd1 vccd1 _6262_/B sky130_fd_sc_hd__clkbuf_2
X_7402_ _7265_/C _7021_/B _7400_/Y _7006_/X vssd1 vssd1 vccd1 vccd1 _7411_/B sky130_fd_sc_hd__a31o_1
X_4614_ _6433_/B vssd1 vssd1 vccd1 vccd1 _5443_/B sky130_fd_sc_hd__clkbuf_2
X_4545_ _7842_/B vssd1 vssd1 vccd1 vccd1 _7943_/B sky130_fd_sc_hd__clkbuf_4
X_7333_ _7333_/A _7333_/B vssd1 vssd1 vccd1 vccd1 _7370_/C sky130_fd_sc_hd__xnor2_1
X_4476_ _4480_/A vssd1 vssd1 vccd1 vccd1 _4476_/Y sky130_fd_sc_hd__inv_2
X_7264_ _6758_/Y _6759_/X _6760_/X vssd1 vssd1 vccd1 vccd1 _7265_/C sky130_fd_sc_hd__a21oi_1
XFILLER_104_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6215_ _6215_/A _6218_/B vssd1 vssd1 vccd1 vccd1 _6294_/B sky130_fd_sc_hd__xnor2_2
X_7195_ _7259_/A _7195_/B vssd1 vssd1 vccd1 vccd1 _7217_/A sky130_fd_sc_hd__xnor2_1
X_6146_ _6144_/A _6228_/A _6153_/B _6145_/Y vssd1 vssd1 vccd1 vccd1 _6224_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_85_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_14 _6460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6077_ _6077_/A _6077_/B vssd1 vssd1 vccd1 vccd1 _6077_/Y sky130_fd_sc_hd__nand2_1
XFILLER_57_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5028_ _5085_/A _5033_/B _5079_/A vssd1 vssd1 vccd1 vccd1 _5042_/D sky130_fd_sc_hd__or3_1
XFILLER_26_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6979_ _7079_/A _7079_/B vssd1 vssd1 vccd1 vccd1 _6980_/A sky130_fd_sc_hd__nand2_1
X_8718_ _8720_/CLK _8718_/D vssd1 vssd1 vccd1 vccd1 _8718_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8649_ _8723_/CLK _8649_/D vssd1 vssd1 vccd1 vccd1 _8649_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6000_ _6000_/A _6000_/B vssd1 vssd1 vccd1 vccd1 _6066_/B sky130_fd_sc_hd__xnor2_1
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8801__18 vssd1 vssd1 vccd1 vccd1 _8801__18/HI _8896_/A sky130_fd_sc_hd__conb_1
XFILLER_67_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7951_ _7951_/A _8022_/B vssd1 vssd1 vccd1 vccd1 _8036_/B sky130_fd_sc_hd__xnor2_1
XFILLER_82_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7882_ _7882_/A _7882_/B vssd1 vssd1 vccd1 vccd1 _8571_/B sky130_fd_sc_hd__xor2_1
X_6902_ _7198_/A _7198_/B vssd1 vssd1 vccd1 vccd1 _7022_/A sky130_fd_sc_hd__nor2_1
X_6833_ _7380_/A vssd1 vssd1 vccd1 vccd1 _7198_/B sky130_fd_sc_hd__buf_2
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6764_ _6764_/A _6764_/B vssd1 vssd1 vccd1 vccd1 _6910_/B sky130_fd_sc_hd__xnor2_4
X_8503_ _8503_/A _8503_/B vssd1 vssd1 vccd1 vccd1 _8544_/A sky130_fd_sc_hd__xnor2_1
X_5715_ _5715_/A vssd1 vssd1 vccd1 vccd1 _5715_/Y sky130_fd_sc_hd__inv_2
X_6695_ _6702_/A _6695_/B vssd1 vssd1 vccd1 vccd1 _6696_/B sky130_fd_sc_hd__nand2_1
X_8434_ _8434_/A vssd1 vssd1 vccd1 vccd1 _8434_/Y sky130_fd_sc_hd__inv_2
X_5646_ _5714_/A _5714_/B vssd1 vssd1 vccd1 vccd1 _5673_/A sky130_fd_sc_hd__xnor2_1
X_8365_ _8284_/A _8284_/B _8364_/Y vssd1 vssd1 vccd1 vccd1 _8435_/A sky130_fd_sc_hd__a21oi_2
X_5577_ _8718_/Q vssd1 vssd1 vccd1 vccd1 _6402_/S sky130_fd_sc_hd__inv_2
X_8296_ _8340_/A _8296_/B vssd1 vssd1 vccd1 vccd1 _8299_/A sky130_fd_sc_hd__xor2_1
X_7316_ _7316_/A _7316_/B vssd1 vssd1 vccd1 vccd1 _7318_/C sky130_fd_sc_hd__xnor2_1
X_4528_ _6742_/B vssd1 vssd1 vccd1 vccd1 _7775_/B sky130_fd_sc_hd__buf_2
X_4459_ _4462_/A vssd1 vssd1 vccd1 vccd1 _4459_/Y sky130_fd_sc_hd__inv_2
X_7247_ _7247_/A _7247_/B vssd1 vssd1 vccd1 vccd1 _7248_/B sky130_fd_sc_hd__and2_1
XFILLER_49_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7178_ _7179_/A _7179_/B vssd1 vssd1 vccd1 vccd1 _7318_/B sky130_fd_sc_hd__nand2_1
X_6129_ _6129_/A _6129_/B vssd1 vssd1 vccd1 vccd1 _6132_/B sky130_fd_sc_hd__xnor2_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8867__84 vssd1 vssd1 vccd1 vccd1 _8867__84/HI _8976_/A sky130_fd_sc_hd__conb_1
XFILLER_5_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5500_ _8709_/Q _6627_/B vssd1 vssd1 vccd1 vccd1 _5500_/X sky130_fd_sc_hd__and2b_1
XFILLER_9_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6480_ _6486_/C _6480_/B _6517_/B vssd1 vssd1 vccd1 vccd1 _6481_/A sky130_fd_sc_hd__and3b_1
X_5431_ _8711_/Q vssd1 vssd1 vccd1 vccd1 _5484_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_99_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8150_ _8086_/A _8086_/B _8149_/X vssd1 vssd1 vccd1 vccd1 _8234_/A sky130_fd_sc_hd__a21oi_4
X_5362_ _5365_/C _5362_/B vssd1 vssd1 vccd1 vccd1 _8687_/D sky130_fd_sc_hd__nor2_1
X_8081_ _8149_/B _8081_/B vssd1 vssd1 vccd1 vccd1 _8086_/A sky130_fd_sc_hd__xnor2_2
X_7101_ _7198_/A _7119_/A vssd1 vssd1 vccd1 vccd1 _7101_/Y sky130_fd_sc_hd__nor2_1
XFILLER_99_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7032_ _7469_/A _7198_/B vssd1 vssd1 vccd1 vccd1 _7038_/A sky130_fd_sc_hd__nor2_1
X_5293_ _4995_/A _5178_/B _5287_/X _5292_/X _4555_/X vssd1 vssd1 vccd1 vccd1 _5293_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8983_ _8983_/A _4479_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[32] sky130_fd_sc_hd__ebufn_8
XFILLER_55_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7934_ _7934_/A _7934_/B _7934_/C _7934_/D vssd1 vssd1 vccd1 vccd1 _7981_/B sky130_fd_sc_hd__nand4_1
XFILLER_70_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7865_ _7866_/A _7866_/B vssd1 vssd1 vccd1 vccd1 _7893_/A sky130_fd_sc_hd__nor2_1
XFILLER_63_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7796_ _7799_/A _7799_/B _7722_/A vssd1 vssd1 vccd1 vccd1 _7912_/B sky130_fd_sc_hd__a21oi_2
X_6816_ _6816_/A _6949_/A _6816_/C vssd1 vssd1 vccd1 vccd1 _6818_/A sky130_fd_sc_hd__nor3_1
XFILLER_11_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6747_ _6764_/A _6764_/B vssd1 vssd1 vccd1 vccd1 _6784_/B sky130_fd_sc_hd__xor2_2
X_6678_ _6678_/A _6678_/B vssd1 vssd1 vccd1 vccd1 _6679_/B sky130_fd_sc_hd__nand2_1
X_8417_ _8417_/A _8417_/B vssd1 vssd1 vccd1 vccd1 _8422_/A sky130_fd_sc_hd__nand2_1
X_5629_ _5632_/A _5979_/B _5979_/C vssd1 vssd1 vccd1 vccd1 _5630_/A sky130_fd_sc_hd__and3_1
X_8348_ _8348_/A _8348_/B vssd1 vssd1 vccd1 vccd1 _8357_/A sky130_fd_sc_hd__nor2_2
X_8279_ _8279_/A _8279_/B _8279_/C vssd1 vssd1 vccd1 vccd1 _8280_/D sky130_fd_sc_hd__nand3_1
XFILLER_78_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5980_ _5980_/A _5994_/B vssd1 vssd1 vccd1 vccd1 _5981_/B sky130_fd_sc_hd__xnor2_2
XFILLER_17_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4931_ _5136_/B _5163_/A vssd1 vssd1 vccd1 vccd1 _5251_/A sky130_fd_sc_hd__or2_1
X_7650_ _7644_/X _7647_/X _7648_/Y _7649_/X _5491_/X vssd1 vssd1 vccd1 vccd1 _8771_/D
+ sky130_fd_sc_hd__o311a_1
X_4862_ _4877_/B _4897_/B _4897_/C _4877_/A vssd1 vssd1 vccd1 vccd1 _5082_/B sky130_fd_sc_hd__or4b_4
XFILLER_60_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6601_ _8754_/Q vssd1 vssd1 vccd1 vccd1 _6851_/A sky130_fd_sc_hd__inv_2
XFILLER_32_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4793_ _4793_/A vssd1 vssd1 vccd1 vccd1 _8666_/D sky130_fd_sc_hd__clkbuf_1
X_7581_ _7578_/Y _7586_/S _7579_/Y _7585_/B vssd1 vssd1 vccd1 vccd1 _7581_/Y sky130_fd_sc_hd__a22oi_1
X_6532_ _8689_/Q _6532_/B _8693_/Q _6532_/D vssd1 vssd1 vccd1 vccd1 _6534_/B sky130_fd_sc_hd__or4_1
X_6463_ _6463_/A vssd1 vssd1 vccd1 vccd1 _8725_/D sky130_fd_sc_hd__clkbuf_1
X_8202_ _8302_/A _8202_/B vssd1 vssd1 vccd1 vccd1 _8204_/B sky130_fd_sc_hd__nor2_1
X_5414_ _8722_/Q vssd1 vssd1 vccd1 vccd1 _6420_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_8133_ _8133_/A _8133_/B vssd1 vssd1 vccd1 vccd1 _8134_/B sky130_fd_sc_hd__xnor2_1
X_6394_ _6394_/A _6394_/B vssd1 vssd1 vccd1 vccd1 _6394_/Y sky130_fd_sc_hd__nand2_1
X_5345_ _8703_/Q _8702_/Q _5344_/X _8704_/Q vssd1 vssd1 vccd1 vccd1 _6562_/A sky130_fd_sc_hd__a31oi_4
XFILLER_99_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8064_ _8165_/C _8172_/B vssd1 vssd1 vccd1 vccd1 _8064_/Y sky130_fd_sc_hd__nor2_1
XFILLER_87_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5276_ _4917_/A _5275_/Y _5199_/B vssd1 vssd1 vccd1 vccd1 _5277_/C sky130_fd_sc_hd__a21oi_1
X_7015_ _7294_/A _7015_/B vssd1 vssd1 vccd1 vccd1 _7016_/B sky130_fd_sc_hd__and2_1
XFILLER_28_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8966_ _8966_/A _4459_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[15] sky130_fd_sc_hd__ebufn_8
XFILLER_15_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7917_ _7917_/A _7925_/A vssd1 vssd1 vccd1 vccd1 _7918_/B sky130_fd_sc_hd__xnor2_1
XFILLER_70_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8897_ _8897_/A _4378_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[16] sky130_fd_sc_hd__ebufn_8
X_7848_ _8025_/A _8349_/A vssd1 vssd1 vccd1 vccd1 _7940_/C sky130_fd_sc_hd__nor2_2
XFILLER_11_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7779_ _7779_/A _7779_/B vssd1 vssd1 vccd1 vccd1 _8349_/A sky130_fd_sc_hd__xnor2_4
XFILLER_23_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8837__54 vssd1 vssd1 vccd1 vccd1 _8837__54/HI _8946_/A sky130_fd_sc_hd__conb_1
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5130_ _5130_/A _5224_/C _5130_/C _5129_/X vssd1 vssd1 vccd1 vccd1 _5130_/X sky130_fd_sc_hd__or4b_1
X_5061_ _5274_/B _5174_/B _5036_/B _5288_/A vssd1 vssd1 vccd1 vccd1 _5064_/C sky130_fd_sc_hd__o31a_1
XFILLER_77_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5963_ _6370_/A _5965_/C _5965_/A vssd1 vssd1 vccd1 vccd1 _6369_/C sky130_fd_sc_hd__o21ai_2
X_8751_ _8753_/CLK _8751_/D vssd1 vssd1 vccd1 vccd1 _8751_/Q sky130_fd_sc_hd__dfxtp_1
X_7702_ _7702_/A _7702_/B vssd1 vssd1 vccd1 vccd1 _8190_/A sky130_fd_sc_hd__xnor2_4
X_4914_ _5189_/B _5135_/B vssd1 vssd1 vccd1 vccd1 _5281_/B sky130_fd_sc_hd__or2_2
X_5894_ _5637_/A _5892_/Y _5893_/X vssd1 vssd1 vccd1 vccd1 _5895_/B sky130_fd_sc_hd__a21oi_1
X_8682_ _8776_/CLK _8682_/D vssd1 vssd1 vccd1 vccd1 _8682_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7633_ _7631_/Y _7633_/B vssd1 vssd1 vccd1 vccd1 _7634_/B sky130_fd_sc_hd__and2b_1
X_4845_ _5007_/A _5157_/B vssd1 vssd1 vccd1 vccd1 _5078_/B sky130_fd_sc_hd__or2_1
X_4776_ _7642_/A vssd1 vssd1 vccd1 vccd1 _7606_/A sky130_fd_sc_hd__buf_2
XFILLER_20_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7564_ _7556_/A _7578_/B _7557_/Y vssd1 vssd1 vccd1 vccd1 _7565_/B sky130_fd_sc_hd__a21o_1
X_6515_ _8742_/Q _6515_/B _6515_/C vssd1 vssd1 vccd1 vccd1 _6519_/B sky130_fd_sc_hd__and3_1
X_7495_ _7419_/A _7419_/B _7494_/Y vssd1 vssd1 vccd1 vccd1 _7498_/A sky130_fd_sc_hd__a21bo_1
X_6446_ _8738_/Q vssd1 vssd1 vccd1 vccd1 _6506_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6377_ _6377_/A _6377_/B vssd1 vssd1 vccd1 vccd1 _6377_/X sky130_fd_sc_hd__or2_1
X_8116_ _8116_/A _8116_/B vssd1 vssd1 vccd1 vccd1 _8117_/B sky130_fd_sc_hd__xnor2_1
X_5328_ _8680_/Q _5334_/B vssd1 vssd1 vccd1 vccd1 _5328_/X sky130_fd_sc_hd__or2_1
XFILLER_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8047_ _8057_/A _8047_/B _8047_/C vssd1 vssd1 vccd1 vccd1 _8057_/B sky130_fd_sc_hd__nand3_1
XFILLER_87_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5259_ _4555_/X _5148_/X _5259_/C _5259_/D vssd1 vssd1 vccd1 vccd1 _5259_/X sky130_fd_sc_hd__and4bb_1
XFILLER_56_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8949_ _8949_/A _4447_/Y vssd1 vssd1 vccd1 vccd1 io_out[36] sky130_fd_sc_hd__ebufn_8
XFILLER_71_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4630_ _4630_/A _4630_/B vssd1 vssd1 vccd1 vccd1 _8634_/D sky130_fd_sc_hd__nor2_1
XFILLER_8_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6300_ _6300_/A _6300_/B vssd1 vssd1 vccd1 vccd1 _6300_/Y sky130_fd_sc_hd__nand2_1
XFILLER_8_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4561_ _5188_/A vssd1 vssd1 vccd1 vccd1 _5066_/A sky130_fd_sc_hd__clkbuf_2
X_4492_ _8656_/Q vssd1 vssd1 vccd1 vccd1 _7729_/B sky130_fd_sc_hd__buf_4
XFILLER_6_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7280_ _7009_/S _6863_/C _7280_/S vssd1 vssd1 vccd1 vccd1 _7281_/B sky130_fd_sc_hd__mux2_1
X_6231_ _6231_/A _6309_/B vssd1 vssd1 vccd1 vccd1 _6232_/B sky130_fd_sc_hd__xnor2_1
XFILLER_103_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6162_ _6162_/A _6162_/B vssd1 vssd1 vccd1 vccd1 _6213_/A sky130_fd_sc_hd__xor2_1
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5113_ _5192_/B _5288_/B _5228_/B vssd1 vssd1 vccd1 vccd1 _5119_/B sky130_fd_sc_hd__or3_1
XFILLER_97_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6093_ _6093_/A _6093_/B vssd1 vssd1 vccd1 vccd1 _6277_/B sky130_fd_sc_hd__nor2_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5044_ _5238_/C _5043_/X _5210_/A vssd1 vssd1 vccd1 vccd1 _5044_/X sky130_fd_sc_hd__o21a_1
XFILLER_38_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6995_ _6820_/A _6820_/B _6953_/B _6994_/Y vssd1 vssd1 vccd1 vccd1 _7063_/A sky130_fd_sc_hd__o31ai_2
X_5946_ _5946_/A _5946_/B _5946_/C vssd1 vssd1 vccd1 vccd1 _6121_/A sky130_fd_sc_hd__and3_1
XFILLER_80_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8734_ _8742_/CLK _8734_/D vssd1 vssd1 vccd1 vccd1 _8734_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5877_ _5801_/A _5803_/A _5885_/B _5876_/X vssd1 vssd1 vccd1 vccd1 _5883_/A sky130_fd_sc_hd__o211a_1
X_8665_ _8776_/CLK _8665_/D vssd1 vssd1 vccd1 vccd1 _8665_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7616_ _7775_/A _7613_/X _7654_/A _7943_/A vssd1 vssd1 vccd1 vccd1 _7616_/X sky130_fd_sc_hd__a31o_1
X_4828_ _4902_/B _4828_/B vssd1 vssd1 vccd1 vccd1 _5298_/C sky130_fd_sc_hd__nand2b_2
X_8596_ _8603_/A _8596_/B vssd1 vssd1 vccd1 vccd1 _8596_/X sky130_fd_sc_hd__or2_1
X_4759_ _4702_/A _4758_/C _4566_/A vssd1 vssd1 vccd1 vccd1 _4760_/C sky130_fd_sc_hd__o21a_1
X_7547_ _7548_/A _7548_/B vssd1 vssd1 vccd1 vccd1 _7551_/B sky130_fd_sc_hd__or2_1
X_7478_ _7489_/A _7388_/S _7384_/B _7383_/B vssd1 vssd1 vccd1 vccd1 _7479_/B sky130_fd_sc_hd__a31o_1
X_6429_ _6429_/A _6429_/B vssd1 vssd1 vccd1 vccd1 _6429_/Y sky130_fd_sc_hd__xnor2_1
X_8807__24 vssd1 vssd1 vccd1 vccd1 _8807__24/HI _8902_/A sky130_fd_sc_hd__conb_1
XFILLER_75_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5800_ _5879_/A _5800_/B vssd1 vssd1 vccd1 vccd1 _5801_/C sky130_fd_sc_hd__nand2_1
XFILLER_50_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6780_ _6780_/A vssd1 vssd1 vccd1 vccd1 _7020_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_35_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5731_ _5730_/B _5730_/C _5730_/A vssd1 vssd1 vccd1 vccd1 _5744_/B sky130_fd_sc_hd__a21o_1
X_8450_ _8450_/A _8450_/B _8165_/B vssd1 vssd1 vccd1 vccd1 _8450_/X sky130_fd_sc_hd__or3b_1
X_5662_ _5916_/A _5662_/B vssd1 vssd1 vccd1 vccd1 _5662_/X sky130_fd_sc_hd__or2_1
XFILLER_30_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8381_ _8381_/A _8381_/B vssd1 vssd1 vccd1 vccd1 _8382_/B sky130_fd_sc_hd__nor2_1
X_5593_ _5688_/A _5993_/A vssd1 vssd1 vccd1 vccd1 _5594_/A sky130_fd_sc_hd__nand2_1
X_4613_ _5462_/A _5462_/B vssd1 vssd1 vccd1 vccd1 _6433_/B sky130_fd_sc_hd__nand2_1
XFILLER_30_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7401_ _7021_/B _7400_/Y _7265_/C vssd1 vssd1 vccd1 vccd1 _7411_/A sky130_fd_sc_hd__a21oi_1
X_7332_ _7332_/A _7366_/A vssd1 vssd1 vccd1 vccd1 _7333_/B sky130_fd_sc_hd__xnor2_1
X_4544_ _8671_/Q vssd1 vssd1 vccd1 vccd1 _7842_/B sky130_fd_sc_hd__clkinv_4
X_7263_ _7279_/A _7279_/B _6792_/B _6836_/A vssd1 vssd1 vccd1 vccd1 _7266_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_104_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6214_ _6217_/B _6214_/B vssd1 vssd1 vccd1 vccd1 _6218_/B sky130_fd_sc_hd__xnor2_1
X_4475_ _4481_/A vssd1 vssd1 vccd1 vccd1 _4480_/A sky130_fd_sc_hd__clkbuf_2
X_7194_ _7194_/A _7194_/B vssd1 vssd1 vccd1 vccd1 _7195_/B sky130_fd_sc_hd__xnor2_2
X_6145_ _6169_/B vssd1 vssd1 vccd1 vccd1 _6145_/Y sky130_fd_sc_hd__clkinv_2
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6076_ _6177_/A _6076_/B vssd1 vssd1 vccd1 vccd1 _6102_/A sky130_fd_sc_hd__and2_2
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_15 _5156_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5027_ _4867_/B _5040_/B _5288_/B vssd1 vssd1 vccd1 vccd1 _5079_/A sky130_fd_sc_hd__o21bai_1
XFILLER_54_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8717_ _8785_/CLK _8717_/D vssd1 vssd1 vccd1 vccd1 _8717_/Q sky130_fd_sc_hd__dfxtp_1
X_6978_ _6978_/A _6978_/B vssd1 vssd1 vccd1 vccd1 _7070_/A sky130_fd_sc_hd__xnor2_1
XFILLER_41_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5929_ _6142_/B _5856_/A _6160_/A vssd1 vssd1 vccd1 vccd1 _5946_/B sky130_fd_sc_hd__a21o_1
XFILLER_70_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8648_ _8723_/CLK _8648_/D vssd1 vssd1 vccd1 vccd1 _8648_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8579_ _8588_/A _8776_/Q vssd1 vssd1 vccd1 vccd1 _8579_/Y sky130_fd_sc_hd__nor2_1
XFILLER_5_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8798__15 vssd1 vssd1 vccd1 vccd1 _8798__15/HI _8893_/A sky130_fd_sc_hd__conb_1
XFILLER_67_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7950_ _7955_/A _8023_/B vssd1 vssd1 vccd1 vccd1 _8022_/B sky130_fd_sc_hd__xnor2_1
XFILLER_67_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7881_ _8568_/C _8249_/A vssd1 vssd1 vccd1 vccd1 _8567_/B sky130_fd_sc_hd__nor2_1
X_6901_ _7182_/A _6910_/C vssd1 vssd1 vccd1 vccd1 _7416_/B sky130_fd_sc_hd__xor2_2
X_6832_ _7036_/A vssd1 vssd1 vccd1 vccd1 _7380_/A sky130_fd_sc_hd__buf_2
XFILLER_23_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6763_ _6774_/A vssd1 vssd1 vccd1 vccd1 _6765_/A sky130_fd_sc_hd__clkinv_2
X_8502_ _8428_/A _8428_/B _8427_/B _8427_/A vssd1 vssd1 vccd1 vccd1 _8503_/B sky130_fd_sc_hd__o2bb2a_1
X_5714_ _5714_/A _5714_/B vssd1 vssd1 vccd1 vccd1 _5714_/X sky130_fd_sc_hd__or2_1
XFILLER_50_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6694_ _6694_/A vssd1 vssd1 vccd1 vccd1 _6825_/A sky130_fd_sc_hd__clkbuf_2
X_8433_ _8433_/A _8433_/B vssd1 vssd1 vccd1 vccd1 _8473_/A sky130_fd_sc_hd__xnor2_1
X_5645_ _6263_/A _6378_/D _5645_/C vssd1 vssd1 vccd1 vccd1 _5714_/B sky130_fd_sc_hd__or3_1
XFILLER_31_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8364_ _8364_/A _8364_/B vssd1 vssd1 vccd1 vccd1 _8364_/Y sky130_fd_sc_hd__nor2_1
X_5576_ _5608_/A _5608_/B vssd1 vssd1 vccd1 vccd1 _5979_/A sky130_fd_sc_hd__xor2_2
X_8295_ _8339_/A _8339_/B vssd1 vssd1 vccd1 vccd1 _8296_/B sky130_fd_sc_hd__xor2_1
X_7315_ _7461_/A _7315_/B vssd1 vssd1 vccd1 vccd1 _7316_/B sky130_fd_sc_hd__nor2_1
XFILLER_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4527_ _8670_/Q vssd1 vssd1 vccd1 vccd1 _6742_/B sky130_fd_sc_hd__inv_2
X_4458_ _4462_/A vssd1 vssd1 vccd1 vccd1 _4458_/Y sky130_fd_sc_hd__inv_2
X_7246_ _7247_/A _7247_/B vssd1 vssd1 vccd1 vccd1 _7248_/A sky130_fd_sc_hd__nor2_1
X_7177_ _7177_/A _7177_/B vssd1 vssd1 vccd1 vccd1 _7179_/B sky130_fd_sc_hd__xnor2_1
X_6128_ _6128_/A _6128_/B vssd1 vssd1 vccd1 vccd1 _6132_/A sky130_fd_sc_hd__nand2_1
X_4389_ _4395_/A vssd1 vssd1 vccd1 vccd1 _4394_/A sky130_fd_sc_hd__clkbuf_2
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6059_ _6059_/A _6228_/A vssd1 vssd1 vccd1 vccd1 _6059_/X sky130_fd_sc_hd__or2_1
XFILLER_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5430_ _8712_/Q vssd1 vssd1 vccd1 vccd1 _5478_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5361_ _8687_/Q _5359_/B _5360_/X vssd1 vssd1 vccd1 vccd1 _5362_/B sky130_fd_sc_hd__o21ai_1
X_8080_ _8080_/A _8080_/B vssd1 vssd1 vccd1 vccd1 _8081_/B sky130_fd_sc_hd__xnor2_1
X_7100_ _7100_/A _7100_/B vssd1 vssd1 vccd1 vccd1 _7104_/A sky130_fd_sc_hd__or2_1
X_5292_ _5179_/D _5281_/X _5289_/X _5291_/X vssd1 vssd1 vccd1 vccd1 _5292_/X sky130_fd_sc_hd__o31a_1
X_7031_ _7031_/A vssd1 vssd1 vccd1 vccd1 _7469_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_67_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8982_ _8982_/A _4478_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[31] sky130_fd_sc_hd__ebufn_8
XFILLER_67_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7933_ _7982_/B _7982_/C _7982_/A vssd1 vssd1 vccd1 vccd1 _7934_/D sky130_fd_sc_hd__a21o_1
XFILLER_82_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7864_ _7970_/A _7864_/B vssd1 vssd1 vccd1 vccd1 _7866_/B sky130_fd_sc_hd__nand2_1
XFILLER_23_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7795_ _7804_/A _7795_/B vssd1 vssd1 vccd1 vccd1 _7912_/A sky130_fd_sc_hd__nand2_2
X_6815_ _7034_/B vssd1 vssd1 vccd1 vccd1 _6816_/A sky130_fd_sc_hd__clkinv_2
XFILLER_11_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6746_ _6632_/A _6632_/B _6629_/A vssd1 vssd1 vccd1 vccd1 _6764_/A sky130_fd_sc_hd__a21oi_4
XFILLER_50_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6677_ _8764_/Q _4754_/A vssd1 vssd1 vccd1 vccd1 _6678_/B sky130_fd_sc_hd__or2b_1
X_8416_ _8360_/A _8360_/B _8358_/Y vssd1 vssd1 vccd1 vccd1 _8423_/A sky130_fd_sc_hd__a21oi_1
X_5628_ _5628_/A _5717_/C vssd1 vssd1 vccd1 vccd1 _5640_/A sky130_fd_sc_hd__xnor2_1
X_8347_ _8286_/A _8286_/B _8346_/X vssd1 vssd1 vccd1 vccd1 _8402_/A sky130_fd_sc_hd__a21oi_1
X_5559_ _8722_/Q _6655_/B vssd1 vssd1 vccd1 vccd1 _5615_/A sky130_fd_sc_hd__and2b_1
X_8278_ _8279_/A _8279_/B _8279_/C vssd1 vssd1 vccd1 vccd1 _8280_/C sky130_fd_sc_hd__a21o_1
X_7229_ _7229_/A _7300_/A vssd1 vssd1 vccd1 vccd1 _7230_/B sky130_fd_sc_hd__xnor2_2
XFILLER_73_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_3_1_0_wb_clk_i clkbuf_3_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_14_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4930_ _5083_/B _4935_/B vssd1 vssd1 vccd1 vccd1 _5163_/A sky130_fd_sc_hd__nor2_2
XFILLER_33_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4861_ _4901_/A _4861_/B _5083_/A vssd1 vssd1 vccd1 vccd1 _5053_/B sky130_fd_sc_hd__or3_1
XFILLER_20_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6600_ _6569_/X _6599_/X _6758_/A _5349_/B vssd1 vssd1 vccd1 vccd1 _8753_/D sky130_fd_sc_hd__o2bb2a_1
XFILLER_32_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7580_ _7583_/A _8746_/Q vssd1 vssd1 vccd1 vccd1 _7585_/B sky130_fd_sc_hd__or2_1
X_4792_ _7642_/A _4792_/B _4796_/B vssd1 vssd1 vccd1 vccd1 _4793_/A sky130_fd_sc_hd__and3_1
X_6531_ _8687_/Q _8686_/Q vssd1 vssd1 vccd1 vccd1 _6534_/A sky130_fd_sc_hd__nand2_1
XFILLER_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6462_ _6455_/B _6524_/B vssd1 vssd1 vccd1 vccd1 _6463_/A sky130_fd_sc_hd__and2b_1
X_8201_ _8201_/A _8201_/B vssd1 vssd1 vccd1 vccd1 _8202_/B sky130_fd_sc_hd__nor2_1
X_6393_ _6394_/A _6394_/B vssd1 vssd1 vccd1 vccd1 _6398_/B sky130_fd_sc_hd__or2_1
X_5413_ _8723_/Q vssd1 vssd1 vccd1 vccd1 _6427_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_8132_ _8228_/A _8132_/B vssd1 vssd1 vccd1 vccd1 _8133_/B sky130_fd_sc_hd__and2_1
X_5344_ _8701_/Q _8700_/Q _5344_/C vssd1 vssd1 vccd1 vccd1 _5344_/X sky130_fd_sc_hd__or3_1
XFILLER_99_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8063_ _8063_/A _8063_/B vssd1 vssd1 vccd1 vccd1 _8153_/B sky130_fd_sc_hd__nand2_1
X_5275_ _5275_/A _5275_/B vssd1 vssd1 vccd1 vccd1 _5275_/Y sky130_fd_sc_hd__nor2_1
XFILLER_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7014_ _7014_/A _7014_/B vssd1 vssd1 vccd1 vccd1 _7015_/B sky130_fd_sc_hd__nand2_1
XFILLER_101_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8965_ _8965_/A _4458_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[14] sky130_fd_sc_hd__ebufn_8
XFILLER_83_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7916_ _7916_/A vssd1 vssd1 vccd1 vccd1 _7925_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_8896_ _8896_/A _4376_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[15] sky130_fd_sc_hd__ebufn_8
XFILLER_55_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7847_ _7940_/A _8102_/B vssd1 vssd1 vccd1 vccd1 _7859_/A sky130_fd_sc_hd__nand2_1
XFILLER_23_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7778_ _7778_/A _7778_/B vssd1 vssd1 vccd1 vccd1 _7779_/B sky130_fd_sc_hd__nand2_2
XFILLER_11_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6729_ _6729_/A _6729_/B vssd1 vssd1 vccd1 vccd1 _6729_/X sky130_fd_sc_hd__or2_1
XFILLER_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8852__69 vssd1 vssd1 vccd1 vccd1 _8852__69/HI _8961_/A sky130_fd_sc_hd__conb_1
XFILLER_87_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5060_ _5215_/A vssd1 vssd1 vccd1 vccd1 _5288_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_77_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5962_ _5962_/A _5962_/B vssd1 vssd1 vccd1 vccd1 _6369_/A sky130_fd_sc_hd__nor2_2
X_8750_ _8753_/CLK _8750_/D vssd1 vssd1 vccd1 vccd1 _8750_/Q sky130_fd_sc_hd__dfxtp_1
X_7701_ _7699_/X _7778_/A vssd1 vssd1 vccd1 vccd1 _7702_/B sky130_fd_sc_hd__and2b_1
XFILLER_52_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4913_ _5164_/A _5189_/C vssd1 vssd1 vccd1 vccd1 _5135_/B sky130_fd_sc_hd__or2_2
X_5893_ _5993_/A _5819_/C _5819_/D _5993_/B _5688_/A vssd1 vssd1 vccd1 vccd1 _5893_/X
+ sky130_fd_sc_hd__o32a_1
X_8681_ _8771_/CLK _8681_/D vssd1 vssd1 vccd1 vccd1 _8681_/Q sky130_fd_sc_hd__dfxtp_1
X_7632_ _7672_/A _7632_/B vssd1 vssd1 vccd1 vccd1 _7633_/B sky130_fd_sc_hd__nand2_1
X_4844_ _4784_/A _4982_/A _4935_/B vssd1 vssd1 vccd1 vccd1 _5157_/B sky130_fd_sc_hd__a21oi_4
XFILLER_33_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7563_ _7563_/A _7563_/B vssd1 vssd1 vccd1 vccd1 _7565_/A sky130_fd_sc_hd__nor2_1
X_4775_ _4807_/A vssd1 vssd1 vccd1 vccd1 _7642_/A sky130_fd_sc_hd__clkbuf_2
X_6514_ _6515_/B _6515_/C _6513_/Y vssd1 vssd1 vccd1 vccd1 _8741_/D sky130_fd_sc_hd__a21oi_1
X_7494_ _7494_/A _7494_/B vssd1 vssd1 vccd1 vccd1 _7494_/Y sky130_fd_sc_hd__nand2_1
X_6445_ _8735_/Q _8733_/Q _6443_/X _6444_/X vssd1 vssd1 vccd1 vccd1 _6445_/X sky130_fd_sc_hd__a31o_1
X_6376_ _6377_/A _6377_/B vssd1 vssd1 vccd1 vccd1 _6381_/A sky130_fd_sc_hd__nand2_1
X_8115_ _8115_/A _8115_/B vssd1 vssd1 vccd1 vccd1 _8116_/B sky130_fd_sc_hd__nand2_1
X_5327_ _8778_/Q _5320_/X _5326_/X _5324_/X vssd1 vssd1 vccd1 vccd1 _8679_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8046_ _8056_/A _8056_/B vssd1 vssd1 vccd1 vccd1 _8047_/C sky130_fd_sc_hd__xor2_1
X_5258_ _4558_/X _5253_/Y _5257_/X _4819_/X vssd1 vssd1 vccd1 vccd1 _5258_/X sky130_fd_sc_hd__o211a_1
XFILLER_75_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5189_ _5261_/B _5189_/B _5189_/C vssd1 vssd1 vccd1 vccd1 _5190_/D sky130_fd_sc_hd__or3_1
XFILLER_83_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8948_ _8948_/A _4449_/Y vssd1 vssd1 vccd1 vccd1 io_out[35] sky130_fd_sc_hd__ebufn_8
XFILLER_73_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4560_ _8652_/Q vssd1 vssd1 vccd1 vccd1 _5188_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4491_ _7794_/B vssd1 vssd1 vccd1 vccd1 _4754_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_6_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6230_ _6230_/A _6230_/B vssd1 vssd1 vccd1 vccd1 _6309_/B sky130_fd_sc_hd__xnor2_1
X_6161_ _6161_/A _6219_/B vssd1 vssd1 vccd1 vccd1 _6162_/B sky130_fd_sc_hd__xnor2_1
XFILLER_69_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5112_ _5160_/A _5142_/C _5112_/C _5030_/Y vssd1 vssd1 vccd1 vccd1 _5112_/X sky130_fd_sc_hd__or4b_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6092_ _6092_/A _6200_/B vssd1 vssd1 vccd1 vccd1 _6095_/A sky130_fd_sc_hd__xnor2_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5043_ _5275_/A _4969_/A _5211_/B _5042_/X vssd1 vssd1 vccd1 vccd1 _5043_/X sky130_fd_sc_hd__o31a_1
XFILLER_38_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6994_ _6994_/A _6994_/B vssd1 vssd1 vccd1 vccd1 _6994_/Y sky130_fd_sc_hd__nand2_1
X_5945_ _5922_/A _5862_/A _5944_/Y vssd1 vssd1 vccd1 vccd1 _5946_/C sky130_fd_sc_hd__o21a_1
X_8733_ _8742_/CLK _8733_/D vssd1 vssd1 vccd1 vccd1 _8733_/Q sky130_fd_sc_hd__dfxtp_1
X_5876_ _5885_/A _5875_/B _5875_/C vssd1 vssd1 vccd1 vccd1 _5876_/X sky130_fd_sc_hd__a21o_1
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8664_ _8758_/CLK _8664_/D vssd1 vssd1 vccd1 vccd1 _8664_/Q sky130_fd_sc_hd__dfxtp_1
X_7615_ _8774_/Q vssd1 vssd1 vccd1 vccd1 _7943_/A sky130_fd_sc_hd__clkbuf_2
X_4827_ _7679_/A _4874_/A vssd1 vssd1 vccd1 vccd1 _4828_/B sky130_fd_sc_hd__nand2_1
X_8595_ _8595_/A _8595_/B vssd1 vssd1 vccd1 vccd1 _8596_/B sky130_fd_sc_hd__xnor2_1
XFILLER_21_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4758_ _5301_/A _5300_/A _4758_/C vssd1 vssd1 vccd1 vccd1 _4760_/B sky130_fd_sc_hd__nand3b_1
XFILLER_5_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7546_ _7541_/X _7545_/X _7606_/A _8756_/Q vssd1 vssd1 vccd1 vccd1 _8756_/D sky130_fd_sc_hd__o2bb2a_1
XFILLER_4_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7477_ _7477_/A _7477_/B vssd1 vssd1 vccd1 vccd1 _7479_/A sky130_fd_sc_hd__xnor2_1
X_4689_ _5266_/A vssd1 vssd1 vccd1 vccd1 _5136_/A sky130_fd_sc_hd__clkbuf_2
X_6428_ _6428_/A _6431_/B vssd1 vssd1 vccd1 vccd1 _6429_/B sky130_fd_sc_hd__nor2_1
X_6359_ _6360_/B _6360_/C _6360_/A vssd1 vssd1 vccd1 vccd1 _6359_/Y sky130_fd_sc_hd__a21oi_1
X_8822__39 vssd1 vssd1 vccd1 vccd1 _8822__39/HI _8917_/A sky130_fd_sc_hd__conb_1
X_8029_ _8044_/A _8030_/B _8034_/A vssd1 vssd1 vccd1 vccd1 _8111_/A sky130_fd_sc_hd__o21a_1
XFILLER_29_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5730_ _5730_/A _5730_/B _5730_/C vssd1 vssd1 vccd1 vccd1 _5744_/A sky130_fd_sc_hd__nand3_1
XFILLER_50_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5661_ _5787_/A _5787_/B vssd1 vssd1 vccd1 vccd1 _5667_/A sky130_fd_sc_hd__xor2_1
X_7400_ _7400_/A _7400_/B vssd1 vssd1 vccd1 vccd1 _7400_/Y sky130_fd_sc_hd__nand2_1
X_8380_ _8380_/A _8461_/S vssd1 vssd1 vccd1 vccd1 _8380_/X sky130_fd_sc_hd__or2_1
X_5592_ _5725_/B vssd1 vssd1 vccd1 vccd1 _5993_/A sky130_fd_sc_hd__clkbuf_2
X_4612_ _8639_/Q _4612_/B _4612_/C vssd1 vssd1 vccd1 vccd1 _5462_/B sky130_fd_sc_hd__or3_1
X_7331_ _7331_/A _7331_/B vssd1 vssd1 vccd1 vccd1 _7366_/A sky130_fd_sc_hd__xnor2_2
X_4543_ _4543_/A _4571_/C vssd1 vssd1 vccd1 vccd1 _4543_/Y sky130_fd_sc_hd__nor2_1
X_7262_ _7400_/A _7262_/B vssd1 vssd1 vccd1 vccd1 _7268_/A sky130_fd_sc_hd__nor2_1
XFILLER_104_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6213_ _6213_/A _6213_/B vssd1 vssd1 vccd1 vccd1 _6214_/B sky130_fd_sc_hd__xnor2_1
X_4474_ _4474_/A vssd1 vssd1 vccd1 vccd1 _4474_/Y sky130_fd_sc_hd__inv_2
X_7193_ _7294_/A _7294_/B vssd1 vssd1 vccd1 vccd1 _7194_/B sky130_fd_sc_hd__xor2_2
X_6144_ _6144_/A _6171_/B vssd1 vssd1 vccd1 vccd1 _6153_/B sky130_fd_sc_hd__xor2_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6075_ _6075_/A _6075_/B _6075_/C vssd1 vssd1 vccd1 vccd1 _6076_/B sky130_fd_sc_hd__or3_1
XFILLER_57_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5026_ _5026_/A vssd1 vssd1 vccd1 vccd1 _5033_/B sky130_fd_sc_hd__clkinv_2
XFILLER_53_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6977_ _7075_/A _7075_/B vssd1 vssd1 vccd1 vccd1 _6978_/A sky130_fd_sc_hd__nand2_1
XFILLER_26_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5928_ _6378_/A _5928_/B vssd1 vssd1 vccd1 vccd1 _6160_/A sky130_fd_sc_hd__or2_1
X_8716_ _8785_/CLK _8716_/D vssd1 vssd1 vccd1 vccd1 _8716_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5859_ _5934_/A _5859_/B vssd1 vssd1 vccd1 vccd1 _5936_/B sky130_fd_sc_hd__nor2_1
X_8647_ _8723_/CLK _8647_/D vssd1 vssd1 vccd1 vccd1 _8647_/Q sky130_fd_sc_hd__dfxtp_1
X_8578_ _8578_/A _8578_/B _8582_/B _8578_/D vssd1 vssd1 vccd1 vccd1 _8578_/X sky130_fd_sc_hd__or4_1
X_7529_ _7529_/A _7529_/B vssd1 vssd1 vccd1 vccd1 _7529_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_79_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7880_ _7880_/A _7880_/B vssd1 vssd1 vccd1 vccd1 _8249_/A sky130_fd_sc_hd__nor2_2
X_6900_ _6900_/A vssd1 vssd1 vccd1 vccd1 _6910_/C sky130_fd_sc_hd__buf_2
XFILLER_35_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6831_ _6760_/X _6758_/Y _6759_/X _6752_/A _6798_/A vssd1 vssd1 vccd1 vccd1 _7036_/A
+ sky130_fd_sc_hd__a311o_2
XFILLER_35_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8501_ _8501_/A _8501_/B vssd1 vssd1 vccd1 vccd1 _8503_/A sky130_fd_sc_hd__xnor2_1
XFILLER_50_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6762_ _7123_/A _6866_/D _6835_/A vssd1 vssd1 vccd1 vccd1 _6778_/B sky130_fd_sc_hd__and3_1
X_5713_ _5677_/A _5677_/B _5676_/A vssd1 vssd1 vccd1 vccd1 _5809_/B sky130_fd_sc_hd__o21ai_2
X_6693_ _6814_/A _6693_/B vssd1 vssd1 vccd1 vccd1 _6970_/A sky130_fd_sc_hd__xnor2_1
X_8432_ _8432_/A vssd1 vssd1 vccd1 vccd1 _8433_/B sky130_fd_sc_hd__inv_2
X_5644_ _5725_/A vssd1 vssd1 vccd1 vccd1 _6263_/A sky130_fd_sc_hd__clkbuf_2
X_8363_ _8363_/A _8363_/B vssd1 vssd1 vccd1 vccd1 _8434_/A sky130_fd_sc_hd__xnor2_2
X_5575_ _5585_/A _5585_/B _5587_/B _5574_/X _5572_/A vssd1 vssd1 vccd1 vccd1 _5608_/B
+ sky130_fd_sc_hd__a311o_4
X_7314_ _7314_/A _7314_/B vssd1 vssd1 vccd1 vccd1 _7315_/B sky130_fd_sc_hd__nor2_1
Xclkbuf_4_3_0_wb_clk_i clkbuf_4_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _8753_/CLK
+ sky130_fd_sc_hd__clkbuf_2
X_8294_ _8197_/A _8197_/B _8293_/Y _8194_/B vssd1 vssd1 vccd1 vccd1 _8339_/B sky130_fd_sc_hd__a22o_1
X_4526_ _4804_/A _4804_/B _4870_/A _4543_/A vssd1 vssd1 vccd1 vccd1 _4814_/C sky130_fd_sc_hd__and4_1
X_4457_ _4457_/A vssd1 vssd1 vccd1 vccd1 _4462_/A sky130_fd_sc_hd__clkbuf_2
X_7245_ _7064_/A _7064_/B _7065_/B _7346_/A vssd1 vssd1 vccd1 vccd1 _7247_/B sky130_fd_sc_hd__a22o_1
X_7176_ _7176_/A _7176_/B vssd1 vssd1 vccd1 vccd1 _7177_/B sky130_fd_sc_hd__nor2_1
XFILLER_98_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6127_ _6363_/A _6363_/B vssd1 vssd1 vccd1 vccd1 _6127_/Y sky130_fd_sc_hd__xnor2_1
X_4388_ _4388_/A vssd1 vssd1 vccd1 vccd1 _4388_/Y sky130_fd_sc_hd__inv_2
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6058_ _6058_/A vssd1 vssd1 vccd1 vccd1 _6252_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_65_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5009_ _5100_/A _5100_/B _5009_/C vssd1 vssd1 vccd1 vccd1 _5187_/A sky130_fd_sc_hd__and3_1
XFILLER_45_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8858__75 vssd1 vssd1 vccd1 vccd1 _8858__75/HI _8967_/A sky130_fd_sc_hd__conb_1
X_5360_ _6567_/A vssd1 vssd1 vccd1 vccd1 _5360_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_99_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5291_ _5291_/A _5291_/B _5291_/C _5291_/D vssd1 vssd1 vccd1 vccd1 _5291_/X sky130_fd_sc_hd__or4_1
XFILLER_99_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7030_ _7030_/A _7391_/B vssd1 vssd1 vccd1 vccd1 _7031_/A sky130_fd_sc_hd__or2_1
XFILLER_95_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8981_ _8981_/A _4477_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[30] sky130_fd_sc_hd__ebufn_8
X_7932_ _7982_/A _7982_/B _7982_/C vssd1 vssd1 vccd1 vccd1 _7934_/C sky130_fd_sc_hd__nand3_1
XFILLER_27_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7863_ _7863_/A _7863_/B vssd1 vssd1 vccd1 vccd1 _7864_/B sky130_fd_sc_hd__nand2_1
XFILLER_35_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7794_ _7794_/A _7794_/B vssd1 vssd1 vccd1 vccd1 _7795_/B sky130_fd_sc_hd__nand2_1
X_6814_ _6814_/A _6814_/B vssd1 vssd1 vccd1 vccd1 _6820_/A sky130_fd_sc_hd__xnor2_1
X_6745_ _6898_/A _7279_/B vssd1 vssd1 vccd1 vccd1 _6786_/A sky130_fd_sc_hd__nor2_2
XFILLER_50_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8415_ _8335_/A _8335_/B _8414_/X vssd1 vssd1 vccd1 vccd1 _8424_/A sky130_fd_sc_hd__a21o_1
X_6676_ _6696_/A _6702_/A _6695_/B _6657_/A vssd1 vssd1 vccd1 vccd1 _6679_/A sky130_fd_sc_hd__a31o_1
X_5627_ _5627_/A _5627_/B vssd1 vssd1 vccd1 vccd1 _5717_/C sky130_fd_sc_hd__xor2_1
X_8346_ _8285_/A _8346_/B vssd1 vssd1 vccd1 vccd1 _8346_/X sky130_fd_sc_hd__and2b_1
X_5558_ _5558_/A _5558_/B vssd1 vssd1 vccd1 vccd1 _5678_/A sky130_fd_sc_hd__xnor2_1
X_4509_ _4509_/A vssd1 vssd1 vccd1 vccd1 _8924_/A sky130_fd_sc_hd__clkbuf_1
X_8277_ _8277_/A _8277_/B vssd1 vssd1 vccd1 vccd1 _8279_/C sky130_fd_sc_hd__xnor2_1
X_7228_ _7228_/A _7228_/B vssd1 vssd1 vccd1 vccd1 _7336_/A sky130_fd_sc_hd__and2_1
X_5489_ _5489_/A vssd1 vssd1 vccd1 vccd1 _8713_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7159_ _7485_/A vssd1 vssd1 vccd1 vccd1 _7332_/A sky130_fd_sc_hd__inv_2
XFILLER_100_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4860_ _4934_/A vssd1 vssd1 vccd1 vccd1 _5083_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_82_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6530_ _8701_/Q _8700_/Q _6529_/X vssd1 vssd1 vccd1 vccd1 _6535_/C sky130_fd_sc_hd__or3b_1
X_4791_ _4791_/A _5040_/A _4543_/A vssd1 vssd1 vccd1 vccd1 _4796_/B sky130_fd_sc_hd__or3b_1
X_6461_ _6508_/B vssd1 vssd1 vccd1 vccd1 _6524_/B sky130_fd_sc_hd__clkbuf_2
X_8200_ _8201_/A _8201_/B vssd1 vssd1 vccd1 vccd1 _8302_/A sky130_fd_sc_hd__and2_1
X_6392_ _6387_/X _6383_/X _6390_/X _6391_/Y vssd1 vssd1 vccd1 vccd1 _8715_/D sky130_fd_sc_hd__a31oi_1
X_5412_ _5411_/Y _5409_/C _5349_/B vssd1 vssd1 vccd1 vccd1 _8703_/D sky130_fd_sc_hd__a21oi_1
X_8131_ _8131_/A _8131_/B vssd1 vssd1 vccd1 vccd1 _8132_/B sky130_fd_sc_hd__nand2_1
X_5343_ _8697_/Q _5342_/X _8699_/Q _8698_/Q vssd1 vssd1 vccd1 vccd1 _5344_/C sky130_fd_sc_hd__o211a_1
XFILLER_99_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8062_ _8376_/A vssd1 vssd1 vccd1 vccd1 _8182_/B sky130_fd_sc_hd__buf_2
X_5274_ _5274_/A _5274_/B _5273_/Y vssd1 vssd1 vccd1 vccd1 _5274_/X sky130_fd_sc_hd__or3b_1
X_7013_ _7014_/A _7014_/B vssd1 vssd1 vccd1 vccd1 _7294_/A sky130_fd_sc_hd__or2_2
XFILLER_101_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8964_ _8964_/A _4456_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[13] sky130_fd_sc_hd__ebufn_8
XFILLER_55_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7915_ _7915_/A _8006_/B vssd1 vssd1 vccd1 vccd1 _7916_/A sky130_fd_sc_hd__or2_1
X_8895_ _8895_/A _4375_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[14] sky130_fd_sc_hd__ebufn_8
X_7846_ _8088_/B vssd1 vssd1 vccd1 vccd1 _8102_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_62_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7777_ _7688_/A _7688_/B _7686_/B _7699_/X _7684_/X vssd1 vssd1 vccd1 vccd1 _7778_/B
+ sky130_fd_sc_hd__a311o_1
XFILLER_23_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4989_ _4563_/X _4985_/Y _4987_/X _4988_/Y _4697_/B vssd1 vssd1 vccd1 vccd1 _4989_/X
+ sky130_fd_sc_hd__o221a_1
X_6728_ _6729_/A _6729_/B vssd1 vssd1 vccd1 vccd1 _6728_/Y sky130_fd_sc_hd__nand2_1
X_6659_ _6660_/A _6660_/B vssd1 vssd1 vccd1 vccd1 _6702_/A sky130_fd_sc_hd__or2_1
X_8329_ _8327_/A _8418_/A _8352_/A _8328_/Y vssd1 vssd1 vccd1 vccd1 _8414_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_3_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8828__45 vssd1 vssd1 vccd1 vccd1 _8828__45/HI _8923_/A sky130_fd_sc_hd__conb_1
XFILLER_2_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5961_ _5965_/A _5961_/B _5965_/C vssd1 vssd1 vccd1 vccd1 _6369_/B sky130_fd_sc_hd__or3_2
XFILLER_65_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7700_ _7700_/A _8772_/Q vssd1 vssd1 vccd1 vccd1 _7778_/A sky130_fd_sc_hd__or2b_1
X_8680_ _8771_/CLK _8680_/D vssd1 vssd1 vccd1 vccd1 _8680_/Q sky130_fd_sc_hd__dfxtp_1
X_4912_ _4935_/A _4912_/B vssd1 vssd1 vccd1 vccd1 _5189_/C sky130_fd_sc_hd__nor2_1
X_5892_ _5892_/A _5993_/B vssd1 vssd1 vccd1 vccd1 _5892_/Y sky130_fd_sc_hd__nor2_1
X_7631_ _7672_/A _7632_/B vssd1 vssd1 vccd1 vccd1 _7631_/Y sky130_fd_sc_hd__nor2_1
X_4843_ _4915_/B vssd1 vssd1 vccd1 vccd1 _4982_/A sky130_fd_sc_hd__inv_2
XFILLER_33_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7562_ _7562_/A _7578_/B vssd1 vssd1 vccd1 vccd1 _7563_/B sky130_fd_sc_hd__nor2_1
X_4774_ _4774_/A _4878_/C vssd1 vssd1 vccd1 vccd1 _4877_/C sky130_fd_sc_hd__nand2_1
X_7493_ _7493_/A _7493_/B vssd1 vssd1 vccd1 vccd1 _7499_/A sky130_fd_sc_hd__xnor2_1
X_6513_ _6515_/B _6515_/C _6524_/B vssd1 vssd1 vccd1 vccd1 _6513_/Y sky130_fd_sc_hd__o21ai_1
X_6444_ _8735_/Q _8734_/Q _8736_/Q vssd1 vssd1 vccd1 vccd1 _6444_/X sky130_fd_sc_hd__a21o_1
X_6375_ _6375_/A _6375_/B _6375_/C _6375_/D vssd1 vssd1 vccd1 vccd1 _6390_/B sky130_fd_sc_hd__or4_4
X_8114_ _8114_/A _8114_/B vssd1 vssd1 vccd1 vccd1 _8115_/B sky130_fd_sc_hd__or2_1
X_5326_ _8679_/Q _5326_/B vssd1 vssd1 vccd1 vccd1 _5326_/X sky130_fd_sc_hd__or2_1
XFILLER_0_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8045_ _8128_/A _8044_/Y _8023_/B _7957_/B vssd1 vssd1 vccd1 vccd1 _8056_/B sky130_fd_sc_hd__a2bb2o_1
X_5257_ _5150_/B _5254_/Y _5256_/X vssd1 vssd1 vccd1 vccd1 _5257_/X sky130_fd_sc_hd__a21o_1
XFILLER_68_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5188_ _5188_/A _5188_/B _5188_/C _5188_/D vssd1 vssd1 vccd1 vccd1 _5188_/X sky130_fd_sc_hd__or4_1
X_8947_ _8947_/A _4452_/Y vssd1 vssd1 vccd1 vccd1 io_out[34] sky130_fd_sc_hd__ebufn_8
XFILLER_71_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7829_ _8158_/A _8380_/A vssd1 vssd1 vccd1 vccd1 _8378_/B sky130_fd_sc_hd__nor2_1
XFILLER_51_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4490_ _8660_/Q vssd1 vssd1 vccd1 vccd1 _7794_/B sky130_fd_sc_hd__clkbuf_4
X_6160_ _6160_/A _6160_/B vssd1 vssd1 vccd1 vccd1 _6219_/B sky130_fd_sc_hd__xnor2_1
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5111_ _5036_/A _5036_/B _5110_/X _4715_/B vssd1 vssd1 vccd1 vccd1 _5112_/C sky130_fd_sc_hd__o31a_1
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6091_ _5749_/A _6192_/B _5751_/A _6194_/A vssd1 vssd1 vccd1 vccd1 _6200_/B sky130_fd_sc_hd__o22a_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5042_ _5042_/A _5275_/B _5238_/B _5042_/D vssd1 vssd1 vccd1 vccd1 _5042_/X sky130_fd_sc_hd__or4_1
XFILLER_84_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6993_ _6956_/A _6956_/B _6992_/X vssd1 vssd1 vccd1 vccd1 _7064_/A sky130_fd_sc_hd__a21o_1
X_5944_ _6169_/A vssd1 vssd1 vccd1 vccd1 _5944_/Y sky130_fd_sc_hd__inv_2
X_8732_ _8732_/CLK _8732_/D vssd1 vssd1 vccd1 vccd1 _8732_/Q sky130_fd_sc_hd__dfxtp_1
X_5875_ _5885_/A _5875_/B _5875_/C vssd1 vssd1 vccd1 vccd1 _5885_/B sky130_fd_sc_hd__nand3_1
XFILLER_21_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8663_ _8758_/CLK _8663_/D vssd1 vssd1 vccd1 vccd1 _8663_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8594_ _8594_/A _8594_/B vssd1 vssd1 vccd1 vccd1 _8595_/B sky130_fd_sc_hd__nand2_1
X_7614_ _8772_/Q _7651_/B vssd1 vssd1 vccd1 vccd1 _7654_/A sky130_fd_sc_hd__or2_1
XFILLER_21_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4826_ _7684_/B _4902_/B vssd1 vssd1 vccd1 vccd1 _4927_/B sky130_fd_sc_hd__xnor2_1
X_7545_ _7552_/A _7552_/B _7548_/B _7545_/D vssd1 vssd1 vccd1 vccd1 _7545_/X sky130_fd_sc_hd__or4_1
X_4757_ _4755_/X _4756_/Y _4705_/X vssd1 vssd1 vccd1 vccd1 _8660_/D sky130_fd_sc_hd__o21a_1
XFILLER_4_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7476_ _7417_/A _7497_/A _7501_/A _7268_/A vssd1 vssd1 vccd1 vccd1 _7477_/B sky130_fd_sc_hd__a2bb2o_1
X_4688_ _5275_/A vssd1 vssd1 vccd1 vccd1 _5266_/A sky130_fd_sc_hd__clkbuf_2
X_6427_ _6427_/A _6427_/B vssd1 vssd1 vccd1 vccd1 _6431_/B sky130_fd_sc_hd__nor2_1
X_6358_ _6358_/A _6358_/B _6358_/C vssd1 vssd1 vccd1 vccd1 _6375_/B sky130_fd_sc_hd__and3_1
X_5309_ _8714_/Q _5307_/X _5308_/X _7621_/A vssd1 vssd1 vccd1 vccd1 _8672_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6289_ _6290_/A _6290_/B _6290_/C vssd1 vssd1 vccd1 vccd1 _6304_/A sky130_fd_sc_hd__o21ai_1
XFILLER_88_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8028_ _8028_/A _8428_/A vssd1 vssd1 vccd1 vccd1 _8034_/A sky130_fd_sc_hd__xnor2_2
XFILLER_75_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5660_ _6147_/A _5531_/X _5556_/Y _5532_/A vssd1 vssd1 vccd1 vccd1 _5787_/B sky130_fd_sc_hd__a211o_1
XFILLER_30_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4611_ _4620_/A _4611_/B _4611_/C _4611_/D vssd1 vssd1 vccd1 vccd1 _4612_/C sky130_fd_sc_hd__or4_1
X_5591_ _6378_/C _6262_/A vssd1 vssd1 vccd1 vccd1 _5645_/C sky130_fd_sc_hd__or2_1
X_7330_ _7391_/B _6725_/A _7300_/A _7377_/A vssd1 vssd1 vccd1 vccd1 _7331_/B sky130_fd_sc_hd__o22a_1
X_4542_ _4778_/A _4850_/A _4541_/X vssd1 vssd1 vccd1 vccd1 _4571_/C sky130_fd_sc_hd__o21a_1
X_4473_ _4474_/A vssd1 vssd1 vccd1 vccd1 _4473_/Y sky130_fd_sc_hd__inv_2
X_7261_ _7261_/A vssd1 vssd1 vccd1 vccd1 _7405_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_104_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6212_ _6212_/A _6221_/B vssd1 vssd1 vccd1 vccd1 _6213_/B sky130_fd_sc_hd__xnor2_1
X_7192_ _7192_/A _7192_/B vssd1 vssd1 vccd1 vccd1 _7294_/B sky130_fd_sc_hd__xnor2_2
XFILLER_97_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6143_ _6142_/Y _6377_/A _5928_/B vssd1 vssd1 vccd1 vccd1 _6152_/A sky130_fd_sc_hd__o21ba_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6074_ _6075_/A _6075_/B _6075_/C vssd1 vssd1 vccd1 vccd1 _6177_/A sky130_fd_sc_hd__o21ai_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5025_ _4947_/A _4889_/B _4887_/X vssd1 vssd1 vccd1 vccd1 _5026_/A sky130_fd_sc_hd__o21a_1
XFILLER_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6976_ _6976_/A _6976_/B vssd1 vssd1 vccd1 vccd1 _6978_/B sky130_fd_sc_hd__xor2_1
X_5927_ _6165_/B vssd1 vssd1 vccd1 vccd1 _5928_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_8715_ _8785_/CLK _8715_/D vssd1 vssd1 vccd1 vccd1 _8715_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5858_ _5872_/A _5858_/B _5862_/A vssd1 vssd1 vccd1 vccd1 _5859_/B sky130_fd_sc_hd__nor3_1
X_8646_ _8723_/CLK _8646_/D vssd1 vssd1 vccd1 vccd1 _8646_/Q sky130_fd_sc_hd__dfxtp_1
X_5789_ _5790_/A _5790_/B vssd1 vssd1 vccd1 vccd1 _5884_/A sky130_fd_sc_hd__nor2_1
X_8577_ _8576_/B _8577_/B vssd1 vssd1 vccd1 vccd1 _8578_/D sky130_fd_sc_hd__and2b_1
X_4809_ _6758_/B _4809_/B vssd1 vssd1 vccd1 vccd1 _4810_/C sky130_fd_sc_hd__or2_1
X_7528_ _7156_/Y _7528_/B vssd1 vssd1 vccd1 vccd1 _7529_/B sky130_fd_sc_hd__and2b_1
X_7459_ _7508_/A _7459_/B vssd1 vssd1 vccd1 vccd1 _7472_/A sky130_fd_sc_hd__xor2_1
XFILLER_1_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6830_ _6973_/A _6973_/B vssd1 vssd1 vccd1 vccd1 _6846_/A sky130_fd_sc_hd__nand2_1
XFILLER_47_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6761_ _6758_/Y _6759_/X _6760_/X vssd1 vssd1 vccd1 vccd1 _6835_/A sky130_fd_sc_hd__a21o_1
XFILLER_35_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8500_ _8500_/A _8500_/B vssd1 vssd1 vccd1 vccd1 _8501_/B sky130_fd_sc_hd__xnor2_1
X_5712_ _5712_/A vssd1 vssd1 vccd1 vccd1 _6394_/A sky130_fd_sc_hd__inv_2
XFILLER_62_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6692_ _7147_/A _6682_/Y _6691_/Y vssd1 vssd1 vccd1 vccd1 _6693_/B sky130_fd_sc_hd__a21oi_1
X_8431_ _8289_/B _8343_/B _8430_/Y vssd1 vssd1 vccd1 vccd1 _8432_/A sky130_fd_sc_hd__a21oi_1
X_5643_ _5643_/A _5716_/B vssd1 vssd1 vccd1 vccd1 _5714_/A sky130_fd_sc_hd__xor2_1
XFILLER_31_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8362_ _8362_/A _8362_/B vssd1 vssd1 vccd1 vccd1 _8363_/B sky130_fd_sc_hd__xor2_1
X_5574_ _6415_/A _6660_/B _6615_/B _5573_/Y vssd1 vssd1 vccd1 vccd1 _5574_/X sky130_fd_sc_hd__o211a_1
X_7313_ _7314_/A _7314_/B vssd1 vssd1 vccd1 vccd1 _7461_/A sky130_fd_sc_hd__and2_1
X_4525_ _4823_/A vssd1 vssd1 vccd1 vccd1 _4543_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_8293_ _8293_/A _8358_/A vssd1 vssd1 vccd1 vccd1 _8293_/Y sky130_fd_sc_hd__nor2_1
X_4456_ _4456_/A vssd1 vssd1 vccd1 vccd1 _4456_/Y sky130_fd_sc_hd__inv_2
X_7244_ _7434_/A _7252_/B vssd1 vssd1 vccd1 vccd1 _7247_/A sky130_fd_sc_hd__xnor2_1
X_4387_ _4388_/A vssd1 vssd1 vccd1 vccd1 _4387_/Y sky130_fd_sc_hd__inv_2
X_7175_ _7006_/X _7262_/B _7274_/A _6792_/B vssd1 vssd1 vccd1 vccd1 _7176_/B sky130_fd_sc_hd__a22o_1
X_6126_ _6293_/A _6293_/B vssd1 vssd1 vccd1 vccd1 _6363_/B sky130_fd_sc_hd__xor2_2
XFILLER_85_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6057_ _6057_/A _6250_/A vssd1 vssd1 vccd1 vccd1 _6065_/A sky130_fd_sc_hd__nand2_1
XFILLER_65_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5008_ _5033_/A vssd1 vssd1 vccd1 vccd1 _5283_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_41_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6959_ _6959_/A _6959_/B vssd1 vssd1 vccd1 vccd1 _7079_/B sky130_fd_sc_hd__xnor2_1
X_8629_ _7602_/A _8628_/Y _4615_/A vssd1 vssd1 vccd1 vccd1 _8629_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_14_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5290_ _5265_/C _5124_/D _5185_/D _5174_/C _5163_/C vssd1 vssd1 vccd1 vccd1 _5291_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_99_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8980_ _8980_/A _4476_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[29] sky130_fd_sc_hd__ebufn_8
X_7931_ _7930_/A _7930_/B _7930_/C vssd1 vssd1 vccd1 vccd1 _7982_/C sky130_fd_sc_hd__a21o_1
XFILLER_27_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7862_ _7863_/A _7863_/B vssd1 vssd1 vccd1 vccd1 _7970_/A sky130_fd_sc_hd__or2_1
XFILLER_63_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7793_ _7794_/A _8660_/Q vssd1 vssd1 vccd1 vccd1 _7804_/A sky130_fd_sc_hd__or2_1
X_6813_ _6856_/A _6813_/B vssd1 vssd1 vccd1 vccd1 _6814_/B sky130_fd_sc_hd__xnor2_1
X_6744_ _6770_/A _6770_/B vssd1 vssd1 vccd1 vccd1 _7279_/B sky130_fd_sc_hd__xor2_4
X_6675_ _6674_/A _6674_/B _6678_/A _6674_/D vssd1 vssd1 vccd1 vccd1 _7379_/B sky130_fd_sc_hd__a22oi_4
X_8414_ _8414_/A _8414_/B vssd1 vssd1 vccd1 vccd1 _8414_/X sky130_fd_sc_hd__and2_1
X_5626_ _5626_/A _5750_/C vssd1 vssd1 vccd1 vccd1 _5627_/B sky130_fd_sc_hd__xnor2_1
X_8345_ _8345_/A _8345_/B vssd1 vssd1 vccd1 vccd1 _8403_/A sky130_fd_sc_hd__xor2_1
X_5557_ _5558_/A _5558_/B _5556_/Y _5531_/X vssd1 vssd1 vccd1 vccd1 _5677_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_104_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8276_ _8389_/A _8389_/B vssd1 vssd1 vccd1 vccd1 _8277_/B sky130_fd_sc_hd__or2_1
X_4508_ _4573_/A _4744_/A vssd1 vssd1 vccd1 vccd1 _4509_/A sky130_fd_sc_hd__or2_2
X_5488_ _7589_/A _5488_/B _5488_/C vssd1 vssd1 vccd1 vccd1 _5489_/A sky130_fd_sc_hd__and3_1
X_4439_ _4457_/A vssd1 vssd1 vccd1 vccd1 _4444_/A sky130_fd_sc_hd__buf_2
X_7227_ _7227_/A _7227_/B vssd1 vssd1 vccd1 vccd1 _7235_/A sky130_fd_sc_hd__nand2_1
XFILLER_76_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7158_ _7530_/A _7530_/B _7156_/Y _7157_/Y vssd1 vssd1 vccd1 vccd1 _7525_/C sky130_fd_sc_hd__a211o_1
X_6109_ _6302_/A _6140_/B vssd1 vssd1 vccd1 vccd1 _6110_/B sky130_fd_sc_hd__xor2_1
XFILLER_86_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7089_ _7110_/B _7110_/A vssd1 vssd1 vccd1 vccd1 _7092_/B sky130_fd_sc_hd__or2b_1
XFILLER_58_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4790_ _5334_/B _5040_/A _4543_/A vssd1 vssd1 vccd1 vccd1 _4792_/B sky130_fd_sc_hd__o21bai_1
XFILLER_32_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6460_ _6460_/A _8628_/A vssd1 vssd1 vccd1 vccd1 _6508_/B sky130_fd_sc_hd__and2_2
X_6391_ _8574_/A _8715_/Q vssd1 vssd1 vccd1 vccd1 _6391_/Y sky130_fd_sc_hd__nor2_1
X_5411_ _8703_/Q vssd1 vssd1 vccd1 vccd1 _5411_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8130_ _8131_/A _8131_/B vssd1 vssd1 vccd1 vccd1 _8228_/A sky130_fd_sc_hd__or2_1
X_5342_ _8695_/Q _8694_/Q _5341_/X _8696_/Q vssd1 vssd1 vccd1 vccd1 _5342_/X sky130_fd_sc_hd__a31o_1
X_8061_ _8061_/A _8061_/B vssd1 vssd1 vccd1 vccd1 _8151_/A sky130_fd_sc_hd__nand2_1
XFILLER_87_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5273_ _5145_/B _5087_/B _5033_/B _5272_/X vssd1 vssd1 vccd1 vccd1 _5273_/Y sky130_fd_sc_hd__o31ai_1
X_7012_ _7412_/A _7261_/A vssd1 vssd1 vccd1 vccd1 _7014_/B sky130_fd_sc_hd__xnor2_1
XFILLER_68_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8963_ _8963_/A _4455_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[12] sky130_fd_sc_hd__ebufn_8
X_7914_ _7804_/A _7807_/B _7809_/A _8381_/A vssd1 vssd1 vccd1 vccd1 _8006_/B sky130_fd_sc_hd__a31o_1
X_8894_ _8894_/A _4374_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[13] sky130_fd_sc_hd__ebufn_8
XFILLER_24_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7845_ _7845_/A _7845_/B vssd1 vssd1 vccd1 vccd1 _8088_/B sky130_fd_sc_hd__xor2_2
X_7776_ _7776_/A _7775_/Y vssd1 vssd1 vccd1 vccd1 _7779_/A sky130_fd_sc_hd__or2b_2
X_4988_ _5148_/A _5050_/D vssd1 vssd1 vccd1 vccd1 _4988_/Y sky130_fd_sc_hd__nor2_1
XFILLER_23_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6727_ _6691_/B _6724_/Y _6726_/Y vssd1 vssd1 vccd1 vccd1 _6729_/B sky130_fd_sc_hd__o21ai_1
X_6658_ _8762_/Q vssd1 vssd1 vccd1 vccd1 _6660_/A sky130_fd_sc_hd__inv_2
X_5609_ _5725_/A _5993_/A vssd1 vssd1 vccd1 vccd1 _5609_/Y sky130_fd_sc_hd__nand2_1
X_8328_ _8355_/A vssd1 vssd1 vccd1 vccd1 _8328_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6589_ _6584_/B _6586_/B _6582_/Y vssd1 vssd1 vccd1 vccd1 _6590_/C sky130_fd_sc_hd__a21oi_1
X_8259_ _8264_/A _8173_/B _8258_/X vssd1 vssd1 vccd1 vccd1 _8268_/A sky130_fd_sc_hd__a21o_1
XFILLER_78_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5960_ _5881_/B _5881_/C _5881_/A vssd1 vssd1 vccd1 vccd1 _5965_/C sky130_fd_sc_hd__a21oi_1
XFILLER_37_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5891_ _5891_/A _5993_/B vssd1 vssd1 vccd1 vccd1 _6183_/B sky130_fd_sc_hd__or2_2
XFILLER_52_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4911_ _4934_/B _4926_/B vssd1 vssd1 vccd1 vccd1 _5164_/A sky130_fd_sc_hd__nor2_1
X_7630_ _7630_/A _8767_/Q vssd1 vssd1 vccd1 vccd1 _7632_/B sky130_fd_sc_hd__xor2_1
XFILLER_33_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4842_ _4878_/C _8663_/Q _8664_/Q _4878_/A vssd1 vssd1 vccd1 vccd1 _4915_/B sky130_fd_sc_hd__and4b_1
XFILLER_33_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7561_ _7562_/A _7578_/B vssd1 vssd1 vccd1 vccd1 _7563_/A sky130_fd_sc_hd__and2_1
X_4773_ _5315_/A vssd1 vssd1 vccd1 vccd1 _5313_/B sky130_fd_sc_hd__clkbuf_2
X_7492_ _7412_/A _7412_/B _7491_/X vssd1 vssd1 vccd1 vccd1 _7493_/B sky130_fd_sc_hd__a21oi_1
X_6512_ _6515_/C _6512_/B vssd1 vssd1 vccd1 vccd1 _8740_/D sky130_fd_sc_hd__nor2_1
X_6443_ _6482_/A _8730_/Q _6442_/X _8732_/Q vssd1 vssd1 vccd1 vccd1 _6443_/X sky130_fd_sc_hd__a211o_1
X_6374_ _6365_/X _6366_/Y _6373_/Y vssd1 vssd1 vccd1 vccd1 _6375_/D sky130_fd_sc_hd__a21o_1
X_8113_ _8113_/A _8113_/B vssd1 vssd1 vccd1 vccd1 _8115_/A sky130_fd_sc_hd__nand2_1
X_5325_ _8777_/Q _5320_/X _5323_/X _5324_/X vssd1 vssd1 vccd1 vccd1 _8678_/D sky130_fd_sc_hd__o211a_1
XFILLER_87_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8044_ _8044_/A _8044_/B vssd1 vssd1 vccd1 vccd1 _8044_/Y sky130_fd_sc_hd__nor2_1
X_5256_ _4716_/A _5142_/Y _5141_/X _5255_/Y _5259_/C vssd1 vssd1 vccd1 vccd1 _5256_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_68_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5187_ _5187_/A _5261_/D vssd1 vssd1 vccd1 vccd1 _5265_/C sky130_fd_sc_hd__or2_1
XFILLER_28_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8946_ _8946_/A _4454_/Y vssd1 vssd1 vccd1 vccd1 io_out[33] sky130_fd_sc_hd__ebufn_8
XFILLER_56_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7828_ _7902_/B _7828_/B vssd1 vssd1 vccd1 vccd1 _8380_/A sky130_fd_sc_hd__and2_1
X_7759_ _7759_/A _7759_/B vssd1 vssd1 vccd1 vccd1 _7760_/B sky130_fd_sc_hd__nand2_1
XFILLER_11_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6090_ _5988_/A _6088_/Y _6278_/A vssd1 vssd1 vccd1 vccd1 _6190_/A sky130_fd_sc_hd__o21a_1
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5110_ _5225_/B _5153_/C _5197_/A _5127_/A vssd1 vssd1 vccd1 vccd1 _5110_/X sky130_fd_sc_hd__or4_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5041_ _5041_/A vssd1 vssd1 vccd1 vccd1 _5238_/B sky130_fd_sc_hd__clkbuf_2
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
XFILLER_92_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6992_ _6955_/A _6992_/B vssd1 vssd1 vccd1 vccd1 _6992_/X sky130_fd_sc_hd__and2b_1
X_8731_ _8732_/CLK _8731_/D vssd1 vssd1 vccd1 vccd1 _8731_/Q sky130_fd_sc_hd__dfxtp_1
X_5943_ _6107_/B _5943_/B vssd1 vssd1 vccd1 vccd1 _5946_/A sky130_fd_sc_hd__or2_1
XFILLER_53_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5874_ _5884_/A _5884_/B vssd1 vssd1 vccd1 vccd1 _5875_/C sky130_fd_sc_hd__xor2_1
XFILLER_80_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8662_ _8758_/CLK _8662_/D vssd1 vssd1 vccd1 vccd1 _8662_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8593_ _8593_/A _8766_/Q vssd1 vssd1 vccd1 vccd1 _8594_/B sky130_fd_sc_hd__or2b_1
X_7613_ _7630_/A _8768_/Q _7651_/B _7637_/A _7649_/A vssd1 vssd1 vccd1 vccd1 _7613_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_21_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4825_ _7679_/A _4874_/A vssd1 vssd1 vccd1 vccd1 _4902_/B sky130_fd_sc_hd__nor2_1
XFILLER_21_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7544_ _7544_/A _7544_/B vssd1 vssd1 vccd1 vccd1 _7545_/D sky130_fd_sc_hd__and2_1
X_4756_ _5300_/A _4758_/C vssd1 vssd1 vccd1 vccd1 _4756_/Y sky130_fd_sc_hd__nor2_1
X_4687_ _5172_/A vssd1 vssd1 vccd1 vccd1 _5275_/A sky130_fd_sc_hd__clkbuf_2
X_7475_ _6966_/B _7266_/B _7268_/A _7006_/X vssd1 vssd1 vccd1 vccd1 _7477_/A sky130_fd_sc_hd__a211o_1
X_6426_ _6427_/A _6427_/B vssd1 vssd1 vccd1 vccd1 _6428_/A sky130_fd_sc_hd__and2_1
X_6357_ _6358_/A _6358_/B _6358_/C vssd1 vssd1 vccd1 vccd1 _6375_/A sky130_fd_sc_hd__a21oi_1
XFILLER_102_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5308_ _8672_/Q _5313_/B vssd1 vssd1 vccd1 vccd1 _5308_/X sky130_fd_sc_hd__or2_1
XFILLER_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6288_ _6288_/A _6288_/B vssd1 vssd1 vccd1 vccd1 _6290_/C sky130_fd_sc_hd__xor2_1
XFILLER_88_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8027_ _8109_/A vssd1 vssd1 vccd1 vccd1 _8428_/A sky130_fd_sc_hd__buf_2
X_5239_ _5139_/A _5202_/X _5226_/Y _4716_/A vssd1 vssd1 vccd1 vccd1 _5239_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_56_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8929_ _8929_/A _4416_/Y vssd1 vssd1 vccd1 vccd1 io_out[16] sky130_fd_sc_hd__ebufn_8
XFILLER_71_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4610_ _8647_/Q _8650_/Q _8649_/Q vssd1 vssd1 vccd1 vccd1 _4611_/D sky130_fd_sc_hd__or3_1
XFILLER_30_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5590_ _5984_/C vssd1 vssd1 vccd1 vccd1 _6262_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_30_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4541_ _4901_/A vssd1 vssd1 vccd1 vccd1 _4541_/X sky130_fd_sc_hd__clkbuf_2
X_4472_ _4474_/A vssd1 vssd1 vccd1 vccd1 _4472_/Y sky130_fd_sc_hd__inv_2
X_7260_ _7217_/A _7217_/B _7259_/X vssd1 vssd1 vccd1 vccd1 _7354_/B sky130_fd_sc_hd__a21bo_1
X_6211_ _6243_/A _6211_/B vssd1 vssd1 vccd1 vccd1 _6221_/B sky130_fd_sc_hd__xnor2_1
X_7191_ _7272_/A _7191_/B vssd1 vssd1 vccd1 vccd1 _7192_/B sky130_fd_sc_hd__nor2_1
X_6142_ _6147_/A _6142_/B vssd1 vssd1 vccd1 vccd1 _6142_/Y sky130_fd_sc_hd__nor2_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6073_ _6183_/A _6318_/A _6180_/B vssd1 vssd1 vccd1 vccd1 _6075_/C sky130_fd_sc_hd__mux2_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5024_ _5153_/C _5086_/A vssd1 vssd1 vccd1 vccd1 _5211_/A sky130_fd_sc_hd__or2_1
XFILLER_81_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6975_ _6975_/A _6975_/B vssd1 vssd1 vccd1 vccd1 _7075_/B sky130_fd_sc_hd__and2_1
X_5926_ _5926_/A _6312_/S vssd1 vssd1 vccd1 vccd1 _5943_/B sky130_fd_sc_hd__nor2_1
XFILLER_80_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8714_ _8785_/CLK _8714_/D vssd1 vssd1 vccd1 vccd1 _8714_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8645_ _8723_/CLK _8645_/D vssd1 vssd1 vccd1 vccd1 _8645_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5857_ _5872_/A _5858_/B _5862_/A vssd1 vssd1 vccd1 vccd1 _5934_/A sky130_fd_sc_hd__o21a_1
X_5788_ _5667_/A _5667_/B _5787_/Y vssd1 vssd1 vccd1 vccd1 _5790_/B sky130_fd_sc_hd__a21oi_1
X_8576_ _8577_/B _8576_/B vssd1 vssd1 vccd1 vccd1 _8582_/B sky130_fd_sc_hd__and2b_1
X_4808_ _6758_/B _4809_/B vssd1 vssd1 vccd1 vccd1 _4810_/B sky130_fd_sc_hd__nand2_1
X_8879__96 vssd1 vssd1 vccd1 vccd1 _8879__96/HI _8988_/A sky130_fd_sc_hd__conb_1
X_4739_ _4740_/A _4973_/A vssd1 vssd1 vccd1 vccd1 _4741_/A sky130_fd_sc_hd__and2_1
X_7527_ _7530_/A _7530_/B _7157_/Y vssd1 vssd1 vccd1 vccd1 _7529_/A sky130_fd_sc_hd__a21o_1
X_7458_ _7410_/A _7410_/B _7457_/X vssd1 vssd1 vccd1 vccd1 _7459_/B sky130_fd_sc_hd__a21oi_1
X_6409_ _6409_/A _6415_/B vssd1 vssd1 vccd1 vccd1 _6413_/A sky130_fd_sc_hd__xnor2_1
XFILLER_1_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7389_ _7389_/A _7389_/B vssd1 vssd1 vccd1 vccd1 _7390_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6760_ _6760_/A vssd1 vssd1 vccd1 vccd1 _6760_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5711_ _5711_/A _5711_/B vssd1 vssd1 vccd1 vccd1 _5712_/A sky130_fd_sc_hd__and2_1
X_6691_ _6834_/B _6691_/B vssd1 vssd1 vccd1 vccd1 _6691_/Y sky130_fd_sc_hd__nor2_1
XFILLER_31_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8430_ _8341_/A _8341_/B _8342_/A vssd1 vssd1 vccd1 vccd1 _8430_/Y sky130_fd_sc_hd__a21oi_1
X_5642_ _6378_/D _6262_/B _5642_/C vssd1 vssd1 vccd1 vccd1 _5716_/B sky130_fd_sc_hd__and3_1
X_8361_ _8527_/A _8437_/B vssd1 vssd1 vccd1 vccd1 _8362_/B sky130_fd_sc_hd__xnor2_1
X_5573_ _8720_/Q vssd1 vssd1 vccd1 vccd1 _5573_/Y sky130_fd_sc_hd__inv_2
X_7312_ _7469_/A _7312_/B vssd1 vssd1 vccd1 vccd1 _7314_/B sky130_fd_sc_hd__xnor2_1
X_4524_ _6630_/B vssd1 vssd1 vccd1 vccd1 _4823_/A sky130_fd_sc_hd__clkbuf_2
X_8292_ _8505_/A _8292_/B vssd1 vssd1 vccd1 vccd1 _8339_/A sky130_fd_sc_hd__xnor2_1
X_4455_ _4456_/A vssd1 vssd1 vccd1 vccd1 _4455_/Y sky130_fd_sc_hd__inv_2
X_7243_ _7243_/A _7251_/A vssd1 vssd1 vccd1 vccd1 _7252_/B sky130_fd_sc_hd__xnor2_1
XFILLER_98_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4386_ _4388_/A vssd1 vssd1 vccd1 vccd1 _4386_/Y sky130_fd_sc_hd__inv_2
X_7174_ _7280_/S vssd1 vssd1 vccd1 vccd1 _7274_/A sky130_fd_sc_hd__clkbuf_2
X_6125_ _6125_/A _6125_/B vssd1 vssd1 vccd1 vccd1 _6293_/B sky130_fd_sc_hd__xnor2_2
XFILLER_100_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6056_ _6029_/A _6029_/B _6055_/Y vssd1 vssd1 vccd1 vccd1 _6137_/A sky130_fd_sc_hd__a21oi_2
XFILLER_100_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5007_ _5007_/A _5149_/B vssd1 vssd1 vccd1 vccd1 _5188_/C sky130_fd_sc_hd__or2_1
XFILLER_81_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6958_ _6958_/A _7078_/B vssd1 vssd1 vccd1 vccd1 _6959_/A sky130_fd_sc_hd__nand2_1
X_5909_ _5907_/Y _5908_/X _5897_/A vssd1 vssd1 vccd1 vccd1 _6024_/A sky130_fd_sc_hd__a21oi_2
X_6889_ _6889_/A _6889_/B vssd1 vssd1 vccd1 vccd1 _6892_/B sky130_fd_sc_hd__xnor2_1
X_8628_ _8628_/A _8628_/B vssd1 vssd1 vccd1 vccd1 _8628_/Y sky130_fd_sc_hd__nor2_1
XFILLER_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8559_ _8559_/A _8559_/B _8559_/C vssd1 vssd1 vccd1 vccd1 _8561_/A sky130_fd_sc_hd__and3_1
XFILLER_1_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7930_ _7930_/A _7930_/B _7930_/C vssd1 vssd1 vccd1 vccd1 _7982_/B sky130_fd_sc_hd__nand3_1
XFILLER_36_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7861_ _7710_/X _7784_/Y _7959_/B vssd1 vssd1 vccd1 vccd1 _7863_/B sky130_fd_sc_hd__a21bo_1
XFILLER_63_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6812_ _7389_/A vssd1 vssd1 vccd1 vccd1 _6813_/B sky130_fd_sc_hd__buf_2
XFILLER_23_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7792_ _8784_/Q vssd1 vssd1 vccd1 vccd1 _7794_/A sky130_fd_sc_hd__inv_2
XFILLER_51_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6743_ _6757_/B _6755_/A vssd1 vssd1 vccd1 vccd1 _6770_/B sky130_fd_sc_hd__nor2_2
X_6674_ _6674_/A _6674_/B _6678_/A _6674_/D vssd1 vssd1 vccd1 vccd1 _7363_/B sky130_fd_sc_hd__and4_2
XFILLER_50_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8413_ _8362_/A _8362_/B _8363_/B _8363_/A vssd1 vssd1 vccd1 vccd1 _8506_/B sky130_fd_sc_hd__a2bb2o_1
X_5625_ _5625_/A _5625_/B vssd1 vssd1 vccd1 vccd1 _5750_/C sky130_fd_sc_hd__xnor2_1
XFILLER_31_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8344_ _8344_/A _8409_/B vssd1 vssd1 vccd1 vccd1 _8345_/B sky130_fd_sc_hd__xnor2_1
X_8849__66 vssd1 vssd1 vccd1 vccd1 _8849__66/HI _8958_/A sky130_fd_sc_hd__conb_1
X_5556_ _5556_/A _5556_/B vssd1 vssd1 vccd1 vccd1 _5556_/Y sky130_fd_sc_hd__nand2_1
X_8275_ _8382_/A _8390_/B vssd1 vssd1 vccd1 vccd1 _8277_/A sky130_fd_sc_hd__xor2_1
X_5487_ _5443_/B _5486_/C _5648_/A vssd1 vssd1 vccd1 vccd1 _5488_/C sky130_fd_sc_hd__o21ai_1
X_4507_ _5249_/B _4740_/A _6613_/B vssd1 vssd1 vccd1 vccd1 _4744_/A sky130_fd_sc_hd__and3_1
XFILLER_104_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4438_ _4438_/A vssd1 vssd1 vccd1 vccd1 _4438_/Y sky130_fd_sc_hd__inv_2
X_7226_ _7056_/A _7056_/B _7225_/X vssd1 vssd1 vccd1 vccd1 _7236_/A sky130_fd_sc_hd__o21ai_1
XFILLER_104_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4369_ _4369_/A vssd1 vssd1 vccd1 vccd1 _4369_/Y sky130_fd_sc_hd__inv_2
X_7157_ _7157_/A _7157_/B vssd1 vssd1 vccd1 vccd1 _7157_/Y sky130_fd_sc_hd__nor2_1
X_6108_ _6230_/A _6016_/B _6059_/X vssd1 vssd1 vccd1 vccd1 _6140_/B sky130_fd_sc_hd__o21a_1
XFILLER_58_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7088_ _7078_/A _7078_/B _7082_/B _7087_/Y vssd1 vssd1 vccd1 vccd1 _7110_/A sky130_fd_sc_hd__a31o_1
X_6039_ _5946_/A _5946_/C _5946_/B vssd1 vssd1 vccd1 vccd1 _6040_/B sky130_fd_sc_hd__a21boi_1
XFILLER_73_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8863__80 vssd1 vssd1 vccd1 vccd1 _8863__80/HI _8972_/A sky130_fd_sc_hd__conb_1
XFILLER_96_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6390_ _6390_/A _6390_/B _6394_/B _6390_/D vssd1 vssd1 vccd1 vccd1 _6390_/X sky130_fd_sc_hd__or4_1
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5410_ _5410_/A vssd1 vssd1 vccd1 vccd1 _8702_/D sky130_fd_sc_hd__clkbuf_1
X_5341_ _8691_/Q _8690_/Q _5339_/X _6532_/D _8693_/Q vssd1 vssd1 vccd1 vccd1 _5341_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_99_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8060_ _8060_/A _8060_/B vssd1 vssd1 vccd1 vccd1 _8149_/B sky130_fd_sc_hd__nand2_1
XFILLER_99_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5272_ _5288_/A _5272_/B _5272_/C vssd1 vssd1 vccd1 vccd1 _5272_/X sky130_fd_sc_hd__or3_1
X_7011_ _7011_/A _7185_/A vssd1 vssd1 vccd1 vccd1 _7261_/A sky130_fd_sc_hd__xor2_2
XFILLER_101_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8962_ _8962_/A _4453_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[11] sky130_fd_sc_hd__ebufn_8
X_7913_ _7913_/A _8514_/A vssd1 vssd1 vccd1 vccd1 _7918_/A sky130_fd_sc_hd__nor2_1
XFILLER_70_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8893_ _8893_/A _4373_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[12] sky130_fd_sc_hd__ebufn_8
XFILLER_63_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7844_ _7778_/A _7775_/Y _7778_/B _7776_/A vssd1 vssd1 vccd1 vccd1 _7845_/B sky130_fd_sc_hd__a31o_2
X_7775_ _7775_/A _7775_/B vssd1 vssd1 vccd1 vccd1 _7775_/Y sky130_fd_sc_hd__nand2_1
XFILLER_23_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6726_ _6691_/B _6724_/Y _6725_/Y vssd1 vssd1 vccd1 vccd1 _6726_/Y sky130_fd_sc_hd__a21oi_1
X_4987_ _5280_/A _5107_/A _5107_/B _5264_/A vssd1 vssd1 vccd1 vccd1 _4987_/X sky130_fd_sc_hd__a31o_1
X_6657_ _6657_/A _6657_/B vssd1 vssd1 vccd1 vccd1 _6696_/A sky130_fd_sc_hd__nor2_2
X_5608_ _5608_/A _5608_/B vssd1 vssd1 vccd1 vccd1 _5725_/A sky130_fd_sc_hd__xnor2_2
X_6588_ _6593_/A _6588_/B vssd1 vssd1 vccd1 vccd1 _6597_/A sky130_fd_sc_hd__nand2_1
X_8327_ _8327_/A _8355_/B vssd1 vssd1 vccd1 vccd1 _8352_/A sky130_fd_sc_hd__xor2_2
X_5539_ _6378_/B _5528_/Y _5852_/A vssd1 vssd1 vccd1 vccd1 _5558_/B sky130_fd_sc_hd__o21a_1
XFILLER_3_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8258_ _8258_/A _8258_/B vssd1 vssd1 vccd1 vccd1 _8258_/X sky130_fd_sc_hd__and2_1
X_8189_ _8189_/A _8189_/B vssd1 vssd1 vccd1 vccd1 _8204_/A sky130_fd_sc_hd__nor2_1
X_7209_ _7209_/A _7297_/B vssd1 vssd1 vccd1 vccd1 _7214_/A sky130_fd_sc_hd__xnor2_1
XFILLER_86_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8792__9 vssd1 vssd1 vccd1 vccd1 _8792__9/HI _8887_/A sky130_fd_sc_hd__conb_1
XFILLER_59_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5890_ _5890_/A _5890_/B vssd1 vssd1 vccd1 vccd1 _5977_/A sky130_fd_sc_hd__nand2_1
X_4910_ _4910_/A _4910_/B vssd1 vssd1 vccd1 vccd1 _5189_/B sky130_fd_sc_hd__nor2_1
XFILLER_33_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4841_ _5032_/B _4935_/B vssd1 vssd1 vccd1 vccd1 _5007_/A sky130_fd_sc_hd__nor2_2
XFILLER_60_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7560_ _7556_/A _6567_/X _6569_/X _7559_/X vssd1 vssd1 vccd1 vccd1 _8760_/D sky130_fd_sc_hd__a22o_1
X_4772_ _4791_/A vssd1 vssd1 vccd1 vccd1 _5315_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7491_ _7415_/A _7491_/B vssd1 vssd1 vccd1 vccd1 _7491_/X sky130_fd_sc_hd__and2b_1
X_6511_ _8740_/Q _6510_/B _6465_/X vssd1 vssd1 vccd1 vccd1 _6512_/B sky130_fd_sc_hd__o21ai_1
X_6442_ _8727_/Q _8728_/Q _6482_/A _6452_/A vssd1 vssd1 vccd1 vccd1 _6442_/X sky130_fd_sc_hd__o211a_1
X_8819__36 vssd1 vssd1 vccd1 vccd1 _8819__36/HI _8914_/A sky130_fd_sc_hd__conb_1
X_6373_ _6365_/C _6367_/X _6368_/Y _6369_/X _6372_/Y vssd1 vssd1 vccd1 vccd1 _6373_/Y
+ sky130_fd_sc_hd__o221ai_1
X_8112_ _8189_/A _8189_/B vssd1 vssd1 vccd1 vccd1 _8116_/A sky130_fd_sc_hd__xnor2_1
Xclkbuf_3_0_0_wb_clk_i clkbuf_3_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
X_5324_ _5335_/A vssd1 vssd1 vccd1 vccd1 _5324_/X sky130_fd_sc_hd__clkbuf_2
X_8043_ _8044_/A _8044_/B vssd1 vssd1 vccd1 vccd1 _8128_/A sky130_fd_sc_hd__and2_1
X_5255_ _5255_/A _5272_/C vssd1 vssd1 vccd1 vccd1 _5255_/Y sky130_fd_sc_hd__nor2_1
XFILLER_68_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5186_ _5274_/A _5127_/A _5098_/C _5185_/X vssd1 vssd1 vccd1 vccd1 _5186_/X sky130_fd_sc_hd__o31a_1
XFILLER_95_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8945_ _8945_/A _4488_/Y vssd1 vssd1 vccd1 vccd1 io_out[32] sky130_fd_sc_hd__ebufn_8
XFILLER_71_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7827_ _8073_/A vssd1 vssd1 vccd1 vccd1 _8158_/A sky130_fd_sc_hd__clkbuf_2
X_7758_ _7759_/A _7759_/B vssd1 vssd1 vccd1 vccd1 _7867_/A sky130_fd_sc_hd__or2_1
XFILLER_51_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7689_ _7689_/A _7689_/B vssd1 vssd1 vccd1 vccd1 _8092_/A sky130_fd_sc_hd__nor2_1
X_6709_ _6809_/A _7034_/B vssd1 vssd1 vccd1 vccd1 _6714_/A sky130_fd_sc_hd__or2_2
XFILLER_22_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8833__50 vssd1 vssd1 vccd1 vccd1 _8833__50/HI _8942_/A sky130_fd_sc_hd__conb_1
XFILLER_78_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5040_ _5040_/A _5040_/B vssd1 vssd1 vccd1 vccd1 _5275_/B sky130_fd_sc_hd__nor2_2
XFILLER_97_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6991_ _7485_/A vssd1 vssd1 vccd1 vccd1 _7346_/A sky130_fd_sc_hd__clkbuf_2
X_5942_ _5942_/A _5866_/B vssd1 vssd1 vccd1 vccd1 _5953_/A sky130_fd_sc_hd__or2b_1
XFILLER_92_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8730_ _8730_/CLK _8730_/D vssd1 vssd1 vccd1 vccd1 _8730_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5873_ _5950_/A _5872_/Y _5851_/C _5785_/B vssd1 vssd1 vccd1 vccd1 _5884_/B sky130_fd_sc_hd__a2bb2o_1
X_8661_ _8778_/CLK _8661_/D vssd1 vssd1 vccd1 vccd1 _8661_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_21_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8592_ _8766_/Q _8593_/A vssd1 vssd1 vccd1 vccd1 _8594_/A sky130_fd_sc_hd__or2b_1
X_7612_ _8771_/Q vssd1 vssd1 vccd1 vccd1 _7649_/A sky130_fd_sc_hd__clkbuf_2
X_4824_ _4874_/A _4874_/B vssd1 vssd1 vccd1 vccd1 _4927_/A sky130_fd_sc_hd__or2_1
X_4755_ _5300_/A _4758_/C vssd1 vssd1 vccd1 vccd1 _4755_/X sky130_fd_sc_hd__and2_1
X_7543_ _7544_/A _7544_/B vssd1 vssd1 vccd1 vccd1 _7548_/B sky130_fd_sc_hd__nor2_1
X_7474_ _7425_/A _7425_/B _7473_/X vssd1 vssd1 vccd1 vccd1 _7480_/A sky130_fd_sc_hd__o21a_1
X_4686_ _8652_/Q vssd1 vssd1 vccd1 vccd1 _5172_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6425_ _6423_/C _6432_/S vssd1 vssd1 vccd1 vccd1 _6429_/A sky130_fd_sc_hd__and2b_1
X_6356_ _6356_/A _6356_/B vssd1 vssd1 vccd1 vccd1 _6358_/C sky130_fd_sc_hd__xnor2_2
XFILLER_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5307_ _5320_/A vssd1 vssd1 vccd1 vccd1 _5307_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6287_ _6351_/A _6351_/B vssd1 vssd1 vccd1 vccd1 _6288_/B sky130_fd_sc_hd__xnor2_1
X_8026_ _7946_/A _8120_/A _8198_/A vssd1 vssd1 vccd1 vccd1 _8109_/A sky130_fd_sc_hd__mux2_2
X_5238_ _5275_/B _5238_/B _5238_/C _5291_/C vssd1 vssd1 vccd1 vccd1 _5238_/X sky130_fd_sc_hd__or4_1
XFILLER_68_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5169_ _4946_/A _5278_/A _5165_/X _5168_/X _4697_/B vssd1 vssd1 vccd1 vccd1 _5170_/C
+ sky130_fd_sc_hd__o311a_1
XFILLER_68_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8928_ _8928_/A _4415_/Y vssd1 vssd1 vccd1 vccd1 io_out[15] sky130_fd_sc_hd__ebufn_8
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4540_ _4877_/A vssd1 vssd1 vccd1 vccd1 _4901_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4471_ _4474_/A vssd1 vssd1 vccd1 vccd1 _4471_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6210_ _6244_/A _6244_/B vssd1 vssd1 vccd1 vccd1 _6211_/B sky130_fd_sc_hd__xor2_1
X_7190_ _7190_/A _7485_/B vssd1 vssd1 vccd1 vccd1 _7191_/B sky130_fd_sc_hd__nor2_1
X_6141_ _6378_/B _6107_/B _6110_/B _6140_/Y vssd1 vssd1 vccd1 vccd1 _6155_/A sky130_fd_sc_hd__a31o_1
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6072_ _6274_/A _6093_/B _6185_/C vssd1 vssd1 vccd1 vccd1 _6318_/A sky130_fd_sc_hd__o21ba_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5023_ _5040_/B _4883_/B _5088_/B vssd1 vssd1 vccd1 vccd1 _5086_/A sky130_fd_sc_hd__o21ai_2
XFILLER_93_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6974_ _7080_/D _6968_/B _6967_/X vssd1 vssd1 vccd1 vccd1 _6975_/B sky130_fd_sc_hd__o21bai_1
X_5925_ _5925_/A _5925_/B vssd1 vssd1 vccd1 vccd1 _6312_/S sky130_fd_sc_hd__nand2_1
X_8713_ _8765_/CLK _8713_/D vssd1 vssd1 vccd1 vccd1 _8713_/Q sky130_fd_sc_hd__dfxtp_1
X_5856_ _5856_/A _6238_/A vssd1 vssd1 vccd1 vccd1 _5862_/A sky130_fd_sc_hd__xnor2_2
X_8644_ _8723_/CLK _8644_/D vssd1 vssd1 vccd1 vccd1 _8644_/Q sky130_fd_sc_hd__dfxtp_1
X_4807_ _4807_/A vssd1 vssd1 vccd1 vccd1 _7589_/A sky130_fd_sc_hd__buf_2
X_5787_ _5787_/A _5787_/B vssd1 vssd1 vccd1 vccd1 _5787_/Y sky130_fd_sc_hd__nor2_1
X_8575_ _6387_/X _8570_/X _8573_/X _8574_/Y vssd1 vssd1 vccd1 vccd1 _8775_/D sky130_fd_sc_hd__a31oi_1
XFILLER_21_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4738_ _5181_/A _4742_/A _4737_/X _4705_/X vssd1 vssd1 vccd1 vccd1 _8656_/D sky130_fd_sc_hd__o211a_1
X_7526_ _7528_/B _7525_/C _7525_/A vssd1 vssd1 vccd1 vccd1 _7526_/Y sky130_fd_sc_hd__a21oi_1
X_4669_ _8647_/Q _4670_/C _4668_/Y vssd1 vssd1 vccd1 vccd1 _8647_/D sky130_fd_sc_hd__a21oi_1
X_7457_ _7408_/B _7457_/B vssd1 vssd1 vccd1 vccd1 _7457_/X sky130_fd_sc_hd__and2b_1
X_6408_ _6405_/A _5449_/X _5450_/X _6407_/Y vssd1 vssd1 vccd1 vccd1 _8719_/D sky130_fd_sc_hd__a22o_1
X_7388_ _6799_/A _6825_/A _7388_/S vssd1 vssd1 vccd1 vccd1 _7389_/B sky130_fd_sc_hd__mux2_1
XFILLER_88_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6339_ _6339_/A _6339_/B vssd1 vssd1 vccd1 vccd1 _6340_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8009_ _7917_/A _8157_/A _7918_/B _7918_/A vssd1 vssd1 vccd1 vccd1 _8082_/A sky130_fd_sc_hd__a22o_1
X_8803__20 vssd1 vssd1 vccd1 vccd1 _8803__20/HI _8898_/A sky130_fd_sc_hd__conb_1
XFILLER_48_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5710_ _5710_/A _5710_/B vssd1 vssd1 vccd1 vccd1 _5711_/B sky130_fd_sc_hd__or2_1
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6690_ _6809_/A _7050_/A vssd1 vssd1 vccd1 vccd1 _6691_/B sky130_fd_sc_hd__nor2_1
XFILLER_31_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5641_ _5749_/A _6262_/A vssd1 vssd1 vccd1 vccd1 _5642_/C sky130_fd_sc_hd__nand2_1
XFILLER_31_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8360_ _8360_/A _8360_/B vssd1 vssd1 vccd1 vccd1 _8437_/B sky130_fd_sc_hd__xnor2_1
X_5572_ _5572_/A _5572_/B vssd1 vssd1 vccd1 vccd1 _5587_/B sky130_fd_sc_hd__nor2_1
X_8291_ _8487_/A _8323_/B vssd1 vssd1 vccd1 vccd1 _8292_/B sky130_fd_sc_hd__xor2_1
X_4523_ _8666_/Q vssd1 vssd1 vccd1 vccd1 _6630_/B sky130_fd_sc_hd__clkbuf_4
X_7311_ _7035_/A _7034_/B _7311_/S vssd1 vssd1 vccd1 vccd1 _7312_/B sky130_fd_sc_hd__mux2_1
X_7242_ _7242_/A _7242_/B vssd1 vssd1 vccd1 vccd1 _7251_/A sky130_fd_sc_hd__xnor2_1
XFILLER_104_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4454_ _4456_/A vssd1 vssd1 vccd1 vccd1 _4454_/Y sky130_fd_sc_hd__inv_2
X_4385_ _4388_/A vssd1 vssd1 vccd1 vccd1 _4385_/Y sky130_fd_sc_hd__inv_2
X_7173_ _6757_/A _6757_/B _6757_/C _7400_/B _6851_/Y vssd1 vssd1 vccd1 vccd1 _7280_/S
+ sky130_fd_sc_hd__o311a_1
X_6124_ _6134_/A _6134_/B vssd1 vssd1 vccd1 vccd1 _6125_/B sky130_fd_sc_hd__xor2_2
XFILLER_98_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6055_ _6055_/A _6055_/B vssd1 vssd1 vccd1 vccd1 _6055_/Y sky130_fd_sc_hd__nor2_1
XFILLER_85_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5006_ _5215_/A _5159_/B _5054_/B _5149_/B vssd1 vssd1 vccd1 vccd1 _5006_/X sky130_fd_sc_hd__or4_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6957_ _6957_/A _6973_/A vssd1 vssd1 vccd1 vccd1 _7079_/A sky130_fd_sc_hd__xnor2_1
XFILLER_26_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5908_ _5908_/A _5840_/B vssd1 vssd1 vccd1 vccd1 _5908_/X sky130_fd_sc_hd__or2b_1
X_6888_ _6888_/A _6888_/B vssd1 vssd1 vccd1 vccd1 _6889_/B sky130_fd_sc_hd__xnor2_1
X_5839_ _5907_/A _5907_/B vssd1 vssd1 vccd1 vccd1 _5840_/B sky130_fd_sc_hd__xor2_1
X_8627_ _8622_/A _8626_/X _8627_/S vssd1 vssd1 vccd1 vccd1 _8628_/B sky130_fd_sc_hd__mux2_1
X_8558_ _8558_/A _8558_/B vssd1 vssd1 vccd1 vccd1 _8558_/X sky130_fd_sc_hd__xor2_1
X_7509_ _7367_/A _7507_/Y _7508_/Y vssd1 vssd1 vccd1 vccd1 _7510_/B sky130_fd_sc_hd__a21oi_1
X_8489_ _8472_/A _8472_/B _8488_/X vssd1 vssd1 vccd1 vccd1 _8490_/B sky130_fd_sc_hd__a21oi_1
XFILLER_30_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7860_ _7860_/A _7860_/B vssd1 vssd1 vccd1 vccd1 _7863_/A sky130_fd_sc_hd__xnor2_1
X_8794__11 vssd1 vssd1 vccd1 vccd1 _8794__11/HI _8889_/A sky130_fd_sc_hd__conb_1
XFILLER_48_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6811_ _7311_/S vssd1 vssd1 vccd1 vccd1 _7389_/A sky130_fd_sc_hd__buf_2
XFILLER_35_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7791_ _8165_/C vssd1 vssd1 vccd1 vccd1 _8163_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_50_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6742_ _8753_/Q _6742_/B vssd1 vssd1 vccd1 vccd1 _6755_/A sky130_fd_sc_hd__nor2_1
X_6673_ _7587_/A _6673_/B vssd1 vssd1 vccd1 vccd1 _6674_/A sky130_fd_sc_hd__nand2_1
XFILLER_31_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8412_ _8403_/A _8403_/B _8411_/X vssd1 vssd1 vccd1 vccd1 _8539_/A sky130_fd_sc_hd__a21o_1
X_5624_ _5687_/A _5979_/B _5979_/C vssd1 vssd1 vccd1 vccd1 _5625_/B sky130_fd_sc_hd__and3_1
X_8343_ _8343_/A _8343_/B vssd1 vssd1 vccd1 vccd1 _8409_/B sky130_fd_sc_hd__xnor2_1
X_5555_ _5766_/A _5913_/A _5550_/Y vssd1 vssd1 vccd1 vccd1 _5556_/B sky130_fd_sc_hd__a21o_1
X_8274_ _7925_/A _8378_/C _7999_/A vssd1 vssd1 vccd1 vccd1 _8390_/B sky130_fd_sc_hd__a21oi_2
X_4506_ _4754_/A _4506_/B _5301_/A vssd1 vssd1 vccd1 vccd1 _4573_/A sky130_fd_sc_hd__or3b_1
X_5486_ _5648_/A _6433_/B _5486_/C vssd1 vssd1 vccd1 vccd1 _5488_/B sky130_fd_sc_hd__or3_1
X_4437_ _4438_/A vssd1 vssd1 vccd1 vccd1 _4437_/Y sky130_fd_sc_hd__inv_2
X_7225_ _7231_/A _7225_/B vssd1 vssd1 vccd1 vccd1 _7225_/X sky130_fd_sc_hd__or2_1
XFILLER_104_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7156_ _7096_/B _7096_/C _7096_/A vssd1 vssd1 vccd1 vccd1 _7156_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_98_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6107_ _6107_/A _6107_/B vssd1 vssd1 vccd1 vccd1 _6320_/A sky130_fd_sc_hd__nand2_2
XFILLER_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4368_ _4369_/A vssd1 vssd1 vccd1 vccd1 _4368_/Y sky130_fd_sc_hd__inv_2
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7087_ _7087_/A _7087_/B vssd1 vssd1 vccd1 vccd1 _7087_/Y sky130_fd_sc_hd__nor2_1
X_6038_ _6036_/Y _6038_/B vssd1 vssd1 vccd1 vccd1 _6121_/B sky130_fd_sc_hd__and2b_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7989_ _8439_/A _7902_/B _7828_/B _7996_/A _8073_/A vssd1 vssd1 vccd1 vccd1 _7991_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_14_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_2_0_wb_clk_i clkbuf_4_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _8742_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_45_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5340_ _8692_/Q vssd1 vssd1 vccd1 vccd1 _6532_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_99_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5271_ _5271_/A _5271_/B _5271_/C vssd1 vssd1 vccd1 vccd1 _5271_/X sky130_fd_sc_hd__or3_1
X_7010_ _7010_/A vssd1 vssd1 vccd1 vccd1 _7185_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_68_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8961_ _8961_/A _4450_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[10] sky130_fd_sc_hd__ebufn_8
XFILLER_28_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7912_ _7912_/A _7912_/B vssd1 vssd1 vccd1 vccd1 _8514_/A sky130_fd_sc_hd__xnor2_2
XFILLER_55_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8892_ _8892_/A _4372_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[11] sky130_fd_sc_hd__ebufn_8
X_7843_ _8102_/A _7843_/B vssd1 vssd1 vccd1 vccd1 _7845_/A sky130_fd_sc_hd__and2_1
XFILLER_24_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7774_ _8773_/Q _7775_/B vssd1 vssd1 vccd1 vccd1 _7776_/A sky130_fd_sc_hd__nor2_1
X_4986_ _5042_/A vssd1 vssd1 vccd1 vccd1 _5280_/A sky130_fd_sc_hd__buf_2
XFILLER_51_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6725_ _6725_/A _6725_/B vssd1 vssd1 vccd1 vccd1 _6725_/Y sky130_fd_sc_hd__nor2_1
X_6656_ _5249_/A _8763_/Q vssd1 vssd1 vccd1 vccd1 _6657_/B sky130_fd_sc_hd__and2b_1
X_5607_ _5701_/B _5632_/A vssd1 vssd1 vccd1 vccd1 _5626_/A sky130_fd_sc_hd__nand2_1
X_6587_ _6583_/A _6567_/X _6569_/X _6586_/Y vssd1 vssd1 vccd1 vccd1 _8751_/D sky130_fd_sc_hd__a22o_1
X_5538_ _6107_/A vssd1 vssd1 vccd1 vccd1 _6378_/B sky130_fd_sc_hd__buf_2
X_8326_ _8325_/Y _8567_/A _8497_/A vssd1 vssd1 vccd1 vccd1 _8335_/A sky130_fd_sc_hd__o21ba_1
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8257_ _8179_/A _8254_/B _8178_/B _8256_/Y vssd1 vssd1 vccd1 vccd1 _8364_/A sky130_fd_sc_hd__o31a_1
XFILLER_3_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7208_ _7208_/A _7208_/B vssd1 vssd1 vccd1 vccd1 _7297_/B sky130_fd_sc_hd__xor2_1
X_5469_ _5463_/B _5462_/X _5467_/Y _5468_/X _7606_/A vssd1 vssd1 vccd1 vccd1 _8710_/D
+ sky130_fd_sc_hd__o221a_1
X_8188_ _8234_/A _8234_/B vssd1 vssd1 vccd1 vccd1 _8206_/A sky130_fd_sc_hd__xor2_2
XFILLER_59_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7139_ _7139_/A _7119_/X vssd1 vssd1 vccd1 vccd1 _7140_/A sky130_fd_sc_hd__or2b_1
XFILLER_74_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4840_ _4926_/B vssd1 vssd1 vccd1 vccd1 _4935_/B sky130_fd_sc_hd__buf_2
XFILLER_33_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6510_ _8740_/Q _6510_/B vssd1 vssd1 vccd1 vccd1 _6515_/C sky130_fd_sc_hd__and2_1
X_4771_ _4771_/A _4771_/B vssd1 vssd1 vccd1 vccd1 _4791_/A sky130_fd_sc_hd__and2_1
X_7490_ _7405_/A _7449_/B _7489_/Y vssd1 vssd1 vccd1 vccd1 _7493_/A sky130_fd_sc_hd__a21o_1
X_6441_ _8729_/Q vssd1 vssd1 vccd1 vccd1 _6452_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6372_ _6372_/A _6372_/B vssd1 vssd1 vccd1 vccd1 _6372_/Y sky130_fd_sc_hd__xnor2_1
X_8111_ _8111_/A _8111_/B vssd1 vssd1 vccd1 vccd1 _8189_/B sky130_fd_sc_hd__nor2_1
X_5323_ _8678_/Q _5326_/B vssd1 vssd1 vccd1 vccd1 _5323_/X sky130_fd_sc_hd__or2_1
XFILLER_102_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8042_ _8039_/X _8040_/Y _7981_/X _7964_/X vssd1 vssd1 vccd1 vccd1 _8047_/B sky130_fd_sc_hd__a211o_1
X_5254_ _4920_/A _5219_/A _5096_/B _4950_/X vssd1 vssd1 vccd1 vccd1 _5254_/Y sky130_fd_sc_hd__o31ai_1
XFILLER_102_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5185_ _5288_/A _5274_/A _5238_/B _5185_/D vssd1 vssd1 vccd1 vccd1 _5185_/X sky130_fd_sc_hd__or4_1
XFILLER_95_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8944_ _8944_/A _4435_/Y vssd1 vssd1 vccd1 vccd1 io_out[31] sky130_fd_sc_hd__ebufn_8
XFILLER_71_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7826_ _7826_/A vssd1 vssd1 vccd1 vccd1 _8073_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_24_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7757_ _7998_/A _7757_/B vssd1 vssd1 vccd1 vccd1 _7759_/B sky130_fd_sc_hd__xnor2_1
X_4969_ _4969_/A _5272_/C _5219_/A vssd1 vssd1 vccd1 vccd1 _4969_/X sky130_fd_sc_hd__or3_1
X_7688_ _7688_/A _7688_/B _7688_/C vssd1 vssd1 vccd1 vccd1 _7689_/B sky130_fd_sc_hd__and3_1
X_6708_ _7105_/A _7105_/B vssd1 vssd1 vccd1 vccd1 _6958_/A sky130_fd_sc_hd__and2_1
X_6639_ _6810_/A vssd1 vssd1 vccd1 vccd1 _6707_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_98_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8309_ _8480_/A _8480_/B vssd1 vssd1 vccd1 vccd1 _8552_/B sky130_fd_sc_hd__xor2_2
XFILLER_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6990_ _7120_/A _6810_/A _6799_/A _6943_/A vssd1 vssd1 vccd1 vccd1 _7485_/A sky130_fd_sc_hd__o2bb2a_4
XFILLER_38_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5941_ _5969_/B _5941_/B vssd1 vssd1 vccd1 vccd1 _5955_/A sky130_fd_sc_hd__xnor2_1
XFILLER_92_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5872_ _5872_/A _5872_/B vssd1 vssd1 vccd1 vccd1 _5872_/Y sky130_fd_sc_hd__nor2_1
XFILLER_61_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8660_ _8778_/CLK _8660_/D vssd1 vssd1 vccd1 vccd1 _8660_/Q sky130_fd_sc_hd__dfxtp_4
X_8591_ _8595_/A _8609_/A _8590_/Y vssd1 vssd1 vccd1 vccd1 _8779_/D sky130_fd_sc_hd__a21oi_1
XFILLER_33_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4823_ _4823_/A _4850_/C vssd1 vssd1 vccd1 vccd1 _4874_/B sky130_fd_sc_hd__nor2_1
X_7611_ _8770_/Q vssd1 vssd1 vccd1 vccd1 _7637_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4754_ _4754_/A vssd1 vssd1 vccd1 vccd1 _5300_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_21_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7542_ _7535_/X _7541_/X _7606_/A _8755_/Q vssd1 vssd1 vccd1 vccd1 _8755_/D sky130_fd_sc_hd__o2bb2a_1
X_7473_ _7473_/A _7473_/B vssd1 vssd1 vccd1 vccd1 _7473_/X sky130_fd_sc_hd__or2_1
X_4685_ _4685_/A vssd1 vssd1 vccd1 vccd1 _8651_/D sky130_fd_sc_hd__clkbuf_1
X_6424_ _5450_/A _6422_/Y _6432_/S _5449_/A _6420_/B vssd1 vssd1 vccd1 vccd1 _8722_/D
+ sky130_fd_sc_hd__a32o_1
X_6355_ _6355_/A _6355_/B vssd1 vssd1 vccd1 vccd1 _6356_/B sky130_fd_sc_hd__xnor2_1
X_6286_ _6286_/A _6286_/B vssd1 vssd1 vccd1 vccd1 _6351_/B sky130_fd_sc_hd__xor2_1
X_5306_ _5248_/X _5305_/X _5315_/A vssd1 vssd1 vccd1 vccd1 _5320_/A sky130_fd_sc_hd__a21bo_1
XFILLER_102_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8025_ _8025_/A _8348_/B vssd1 vssd1 vccd1 vccd1 _8198_/A sky130_fd_sc_hd__or2_2
X_5237_ _5124_/D _5197_/C _5116_/A vssd1 vssd1 vccd1 vccd1 _5237_/X sky130_fd_sc_hd__o21a_1
XFILLER_102_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5168_ _5168_/A _5168_/B _5261_/D _4885_/Y vssd1 vssd1 vccd1 vccd1 _5168_/X sky130_fd_sc_hd__or4b_1
X_5099_ _5215_/A _5224_/B _5163_/B _5099_/D vssd1 vssd1 vccd1 vccd1 _5099_/X sky130_fd_sc_hd__or4_1
XFILLER_83_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8927_ _8927_/A _4413_/Y vssd1 vssd1 vccd1 vccd1 io_out[14] sky130_fd_sc_hd__ebufn_8
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7809_ _7809_/A vssd1 vssd1 vccd1 vccd1 _7813_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_33_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4470_ _4474_/A vssd1 vssd1 vccd1 vccd1 _4470_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6140_ _6302_/A _6140_/B vssd1 vssd1 vccd1 vccd1 _6140_/Y sky130_fd_sc_hd__nor2_1
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6071_ _6071_/A _6093_/B vssd1 vssd1 vccd1 vccd1 _6185_/C sky130_fd_sc_hd__and2_1
XFILLER_57_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5022_ _5189_/B _5135_/B vssd1 vssd1 vccd1 vccd1 _5088_/B sky130_fd_sc_hd__nor2_1
XFILLER_65_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6973_ _6973_/A _6973_/B vssd1 vssd1 vccd1 vccd1 _7075_/A sky130_fd_sc_hd__xor2_1
X_5924_ _6036_/A _5923_/X vssd1 vssd1 vccd1 vccd1 _6011_/A sky130_fd_sc_hd__or2b_1
X_8712_ _8720_/CLK _8712_/D vssd1 vssd1 vccd1 vccd1 _8712_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5855_ _5932_/A vssd1 vssd1 vccd1 vccd1 _6238_/A sky130_fd_sc_hd__buf_2
X_8643_ _8723_/CLK _8643_/D vssd1 vssd1 vccd1 vccd1 _8643_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4806_ _4806_/A vssd1 vssd1 vccd1 vccd1 _8669_/D sky130_fd_sc_hd__clkbuf_1
X_5786_ _5786_/A _5786_/B vssd1 vssd1 vccd1 vccd1 _5790_/A sky130_fd_sc_hd__xnor2_1
X_8574_ _8574_/A _8775_/Q vssd1 vssd1 vccd1 vccd1 _8574_/Y sky130_fd_sc_hd__nor2_1
Xclkbuf_4_15_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8776_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_21_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4737_ _4745_/A _5130_/A vssd1 vssd1 vccd1 vccd1 _4737_/X sky130_fd_sc_hd__or2_1
X_7525_ _7525_/A _7528_/B _7525_/C vssd1 vssd1 vccd1 vccd1 _7525_/X sky130_fd_sc_hd__and3_1
XFILLER_21_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4668_ _8647_/Q _4670_/C _4679_/A vssd1 vssd1 vccd1 vccd1 _4668_/Y sky130_fd_sc_hd__o21ai_1
X_7456_ _7456_/A _7456_/B vssd1 vssd1 vccd1 vccd1 _7504_/A sky130_fd_sc_hd__xnor2_1
X_6407_ _8718_/Q _6407_/B vssd1 vssd1 vccd1 vccd1 _6407_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_103_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4599_ _8679_/Q _5305_/A vssd1 vssd1 vccd1 vccd1 _4600_/A sky130_fd_sc_hd__and2_1
X_7387_ _7463_/B _7387_/B vssd1 vssd1 vccd1 vccd1 _7395_/A sky130_fd_sc_hd__xnor2_2
X_6338_ _6338_/A _6338_/B vssd1 vssd1 vccd1 vccd1 _6339_/B sky130_fd_sc_hd__xnor2_1
XFILLER_76_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6269_ _6269_/A _6269_/B vssd1 vssd1 vccd1 vccd1 _6271_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8008_ _8008_/A _8371_/A vssd1 vssd1 vccd1 vccd1 _8083_/A sky130_fd_sc_hd__nand2_1
XFILLER_57_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5640_ _5640_/A _5640_/B vssd1 vssd1 vccd1 vccd1 _5643_/A sky130_fd_sc_hd__xnor2_1
X_5571_ _6660_/B _8721_/Q vssd1 vssd1 vccd1 vccd1 _5572_/B sky130_fd_sc_hd__and2b_1
X_8290_ _8420_/A _8194_/B _8239_/X vssd1 vssd1 vccd1 vccd1 _8323_/B sky130_fd_sc_hd__o21a_1
X_7310_ _6886_/A _7309_/B _7390_/A vssd1 vssd1 vccd1 vccd1 _7314_/A sky130_fd_sc_hd__o21a_1
X_4522_ _7679_/A vssd1 vssd1 vccd1 vccd1 _4870_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4453_ _4456_/A vssd1 vssd1 vccd1 vccd1 _4453_/Y sky130_fd_sc_hd__inv_2
X_7241_ _7241_/A _7253_/A vssd1 vssd1 vccd1 vccd1 _7242_/B sky130_fd_sc_hd__xnor2_1
X_4384_ _4388_/A vssd1 vssd1 vccd1 vccd1 _4384_/Y sky130_fd_sc_hd__inv_2
X_7172_ _7412_/A _7417_/A vssd1 vssd1 vccd1 vccd1 _7177_/A sky130_fd_sc_hd__or2_1
X_6123_ _6123_/A _6123_/B vssd1 vssd1 vccd1 vccd1 _6134_/B sky130_fd_sc_hd__xnor2_2
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6054_ _6045_/A _6045_/B _6053_/X vssd1 vssd1 vccd1 vccd1 _6134_/A sky130_fd_sc_hd__a21boi_2
XFILLER_100_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5005_ _5007_/A _5005_/B vssd1 vssd1 vccd1 vccd1 _5054_/B sky130_fd_sc_hd__or2_1
XFILLER_26_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6956_ _6956_/A _6956_/B vssd1 vssd1 vccd1 vccd1 _6988_/B sky130_fd_sc_hd__xnor2_1
XFILLER_41_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5907_ _5907_/A _5907_/B vssd1 vssd1 vccd1 vccd1 _5907_/Y sky130_fd_sc_hd__nand2_1
X_6887_ _6887_/A _6887_/B vssd1 vssd1 vccd1 vccd1 _6888_/B sky130_fd_sc_hd__xnor2_1
X_5838_ _5980_/A _5838_/B vssd1 vssd1 vccd1 vccd1 _5907_/B sky130_fd_sc_hd__xnor2_1
X_8626_ _8626_/A _8626_/B vssd1 vssd1 vccd1 vccd1 _8626_/X sky130_fd_sc_hd__or2_1
XFILLER_22_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5769_ _5769_/A vssd1 vssd1 vccd1 vccd1 _5769_/Y sky130_fd_sc_hd__inv_2
X_8557_ _8559_/A _8559_/C _8559_/B vssd1 vssd1 vccd1 vccd1 _8558_/B sky130_fd_sc_hd__a21bo_1
X_7508_ _7508_/A _7508_/B vssd1 vssd1 vccd1 vccd1 _7508_/Y sky130_fd_sc_hd__nor2_1
X_8488_ _8473_/A _8488_/B vssd1 vssd1 vccd1 vccd1 _8488_/X sky130_fd_sc_hd__and2b_1
X_7439_ _7521_/A _7437_/X _7438_/X vssd1 vssd1 vccd1 vccd1 _7439_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_76_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6810_ _6810_/A _7302_/A vssd1 vssd1 vccd1 vccd1 _7311_/S sky130_fd_sc_hd__nor2_1
X_7790_ _7904_/A _7899_/A vssd1 vssd1 vccd1 vccd1 _8165_/C sky130_fd_sc_hd__nand2_1
XFILLER_16_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6741_ _8753_/Q _6758_/B vssd1 vssd1 vccd1 vccd1 _6757_/B sky130_fd_sc_hd__and2_1
XFILLER_50_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6672_ _6725_/B vssd1 vssd1 vccd1 vccd1 _7147_/A sky130_fd_sc_hd__inv_2
X_8411_ _8402_/A _8411_/B vssd1 vssd1 vccd1 vccd1 _8411_/X sky130_fd_sc_hd__and2b_1
X_5623_ _5634_/A _5634_/C _5634_/B vssd1 vssd1 vccd1 vccd1 _5979_/C sky130_fd_sc_hd__a21o_1
X_8342_ _8342_/A _8342_/B vssd1 vssd1 vccd1 vccd1 _8343_/B sky130_fd_sc_hd__xnor2_1
X_5554_ _5554_/A _5554_/B vssd1 vssd1 vccd1 vccd1 _5913_/A sky130_fd_sc_hd__xnor2_4
X_8273_ _8273_/A _8273_/B vssd1 vssd1 vccd1 vccd1 _8378_/C sky130_fd_sc_hd__or2_1
X_4505_ _6673_/B vssd1 vssd1 vccd1 vccd1 _5301_/A sky130_fd_sc_hd__clkbuf_1
X_5485_ _5480_/C _5484_/X _5485_/S vssd1 vssd1 vccd1 vccd1 _5486_/C sky130_fd_sc_hd__mux2_1
X_4436_ _4438_/A vssd1 vssd1 vccd1 vccd1 _4436_/Y sky130_fd_sc_hd__inv_2
X_7224_ _7041_/A _7041_/B _7223_/X vssd1 vssd1 vccd1 vccd1 _7238_/A sky130_fd_sc_hd__o21ai_1
XFILLER_98_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4367_ _4369_/A vssd1 vssd1 vccd1 vccd1 _4367_/Y sky130_fd_sc_hd__inv_2
X_7155_ _7519_/A _7519_/B _7154_/X vssd1 vssd1 vccd1 vccd1 _7530_/B sky130_fd_sc_hd__a21o_1
XFILLER_98_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6106_ _6238_/A _6106_/B vssd1 vssd1 vccd1 vccd1 _6157_/A sky130_fd_sc_hd__nand2_1
XFILLER_86_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7086_ _7086_/A _7086_/B vssd1 vssd1 vccd1 vccd1 _7110_/B sky130_fd_sc_hd__xor2_1
XFILLER_100_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6037_ _6036_/A _6036_/C _6036_/B vssd1 vssd1 vccd1 vccd1 _6038_/B sky130_fd_sc_hd__o21ai_1
XFILLER_86_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7988_ _7988_/A _8172_/B vssd1 vssd1 vccd1 vccd1 _8068_/A sky130_fd_sc_hd__nor2_2
XFILLER_81_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6939_ _6939_/A _6939_/B vssd1 vssd1 vccd1 vccd1 _6940_/B sky130_fd_sc_hd__xor2_1
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8609_ _8609_/A _8609_/B vssd1 vssd1 vccd1 vccd1 _8609_/Y sky130_fd_sc_hd__nand2_1
XFILLER_10_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5270_ _5278_/B _5261_/X _5263_/X _5268_/X _5291_/B vssd1 vssd1 vccd1 vccd1 _5271_/C
+ sky130_fd_sc_hd__o32a_1
XFILLER_99_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8854__71 vssd1 vssd1 vccd1 vccd1 _8854__71/HI _8963_/A sky130_fd_sc_hd__conb_1
XFILLER_68_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8960_ _8960_/A _4448_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[9] sky130_fd_sc_hd__ebufn_8
XFILLER_95_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7911_ _7910_/B _7910_/C _7910_/A vssd1 vssd1 vccd1 vccd1 _7919_/B sky130_fd_sc_hd__a21o_1
X_8891_ _8891_/A _4369_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[10] sky130_fd_sc_hd__ebufn_8
X_7842_ _7943_/A _7842_/B vssd1 vssd1 vccd1 vccd1 _7843_/B sky130_fd_sc_hd__nand2_1
XFILLER_36_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7773_ _7773_/A _7872_/B _7773_/C vssd1 vssd1 vccd1 vccd1 _7875_/A sky130_fd_sc_hd__nor3_1
X_4985_ _5224_/B _5005_/B _5199_/A vssd1 vssd1 vccd1 vccd1 _4985_/Y sky130_fd_sc_hd__nor3b_1
X_6724_ _7392_/A _6957_/A vssd1 vssd1 vccd1 vccd1 _6724_/Y sky130_fd_sc_hd__nor2_1
X_6655_ _8763_/Q _6655_/B vssd1 vssd1 vccd1 vccd1 _6657_/A sky130_fd_sc_hd__and2b_1
X_5606_ _5727_/B vssd1 vssd1 vccd1 vccd1 _5632_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6586_ _6586_/A _6586_/B vssd1 vssd1 vccd1 vccd1 _6586_/Y sky130_fd_sc_hd__xnor2_1
X_8325_ _8325_/A _8325_/B vssd1 vssd1 vccd1 vccd1 _8325_/Y sky130_fd_sc_hd__nor2_1
X_5537_ _5681_/A _5535_/B _5684_/A vssd1 vssd1 vccd1 vccd1 _5558_/A sky130_fd_sc_hd__a21o_1
X_8256_ _8256_/A _8256_/B vssd1 vssd1 vccd1 vccd1 _8256_/Y sky130_fd_sc_hd__nand2_1
XFILLER_11_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7207_ _7382_/A _7306_/B vssd1 vssd1 vccd1 vccd1 _7208_/B sky130_fd_sc_hd__xnor2_1
X_5468_ _5467_/A _5467_/B _5443_/B vssd1 vssd1 vccd1 vccd1 _5468_/X sky130_fd_sc_hd__a21o_1
X_4419_ _4419_/A vssd1 vssd1 vccd1 vccd1 _4419_/Y sky130_fd_sc_hd__inv_2
X_8187_ _8187_/A _8187_/B vssd1 vssd1 vccd1 vccd1 _8234_/B sky130_fd_sc_hd__xnor2_4
X_5399_ _8699_/Q _5401_/C _5392_/X vssd1 vssd1 vccd1 vccd1 _5400_/B sky130_fd_sc_hd__o21ai_1
XFILLER_101_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7138_ _7138_/A _7138_/B vssd1 vssd1 vccd1 vccd1 _7145_/B sky130_fd_sc_hd__nor2_1
XFILLER_100_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7069_ _7069_/A _7069_/B vssd1 vssd1 vccd1 vccd1 _7096_/A sky130_fd_sc_hd__xnor2_1
XFILLER_74_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4770_ _4774_/A vssd1 vssd1 vccd1 vccd1 _4897_/B sky130_fd_sc_hd__clkbuf_2
X_6440_ _8731_/Q vssd1 vssd1 vccd1 vccd1 _6482_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6371_ _6369_/A _6369_/C _5965_/Y vssd1 vssd1 vccd1 vccd1 _6372_/B sky130_fd_sc_hd__a21oi_1
XFILLER_9_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8110_ _8110_/A _8487_/A vssd1 vssd1 vccd1 vccd1 _8111_/B sky130_fd_sc_hd__xnor2_1
X_5322_ _8776_/Q _5320_/X _5321_/X _5311_/X vssd1 vssd1 vccd1 vccd1 _8677_/D sky130_fd_sc_hd__o211a_1
X_8041_ _7981_/X _7964_/X _8039_/X _8040_/Y vssd1 vssd1 vccd1 vccd1 _8057_/A sky130_fd_sc_hd__o211ai_2
X_5253_ _5250_/X _5252_/X _5136_/C vssd1 vssd1 vccd1 vccd1 _5253_/Y sky130_fd_sc_hd__a21oi_1
X_5184_ _5189_/B _5184_/B vssd1 vssd1 vccd1 vccd1 _5185_/D sky130_fd_sc_hd__or2_1
XFILLER_3_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8943_ _8943_/A _4434_/Y vssd1 vssd1 vccd1 vccd1 io_out[30] sky130_fd_sc_hd__ebufn_8
X_7825_ _8382_/A vssd1 vssd1 vccd1 vccd1 _7934_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_51_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7756_ _8568_/D _7836_/C _7755_/X vssd1 vssd1 vccd1 vccd1 _7757_/B sky130_fd_sc_hd__o21a_1
X_4968_ _5210_/A _5209_/A vssd1 vssd1 vccd1 vccd1 _5219_/A sky130_fd_sc_hd__or2_1
X_7687_ _7688_/A _7688_/B _7688_/C vssd1 vssd1 vccd1 vccd1 _7689_/A sky130_fd_sc_hd__a21oi_2
X_4899_ _5087_/B _5074_/B vssd1 vssd1 vccd1 vccd1 _5288_/B sky130_fd_sc_hd__or2_2
X_6707_ _6707_/A _7120_/B vssd1 vssd1 vccd1 vccd1 _7105_/B sky130_fd_sc_hd__nor2_1
X_6638_ _6671_/B vssd1 vssd1 vccd1 vccd1 _6810_/A sky130_fd_sc_hd__clkbuf_2
X_8308_ _8308_/A _8308_/B vssd1 vssd1 vccd1 vccd1 _8480_/B sky130_fd_sc_hd__xnor2_2
XFILLER_3_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6569_ _6569_/A vssd1 vssd1 vccd1 vccd1 _6569_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_79_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8239_ _8239_/A _8355_/B vssd1 vssd1 vccd1 vccd1 _8239_/X sky130_fd_sc_hd__or2_1
XFILLER_78_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8824__41 vssd1 vssd1 vccd1 vccd1 _8824__41/HI _8919_/A sky130_fd_sc_hd__conb_1
XFILLER_88_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5940_ _5940_/A _5940_/B vssd1 vssd1 vccd1 vccd1 _5941_/B sky130_fd_sc_hd__xnor2_1
XFILLER_92_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5871_ _5872_/A _5872_/B vssd1 vssd1 vccd1 vccd1 _5950_/A sky130_fd_sc_hd__and2_1
X_7610_ _7637_/B vssd1 vssd1 vccd1 vccd1 _7651_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_8590_ _8595_/A _7649_/B _4615_/A vssd1 vssd1 vccd1 vccd1 _8590_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_21_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4822_ _6630_/B _4850_/C vssd1 vssd1 vccd1 vccd1 _4874_/A sky130_fd_sc_hd__and2_1
X_4753_ _4753_/A vssd1 vssd1 vccd1 vccd1 _8659_/D sky130_fd_sc_hd__clkbuf_1
X_7541_ _7552_/A _7540_/X _7576_/B vssd1 vssd1 vccd1 vccd1 _7541_/X sky130_fd_sc_hd__o21a_1
X_7472_ _7472_/A _7472_/B vssd1 vssd1 vccd1 vccd1 _7481_/A sky130_fd_sc_hd__xnor2_1
X_4684_ _8588_/A _4684_/B vssd1 vssd1 vccd1 vccd1 _4685_/A sky130_fd_sc_hd__and2_1
X_6423_ _6423_/A _6423_/B _6423_/C _6423_/D vssd1 vssd1 vccd1 vccd1 _6432_/S sky130_fd_sc_hd__or4_2
X_6354_ _6354_/A _6354_/B vssd1 vssd1 vccd1 vccd1 _6355_/B sky130_fd_sc_hd__xnor2_1
X_6285_ _6300_/A _6300_/B vssd1 vssd1 vccd1 vccd1 _6286_/B sky130_fd_sc_hd__xor2_1
XFILLER_88_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5305_ _5305_/A _5305_/B _5305_/C _5305_/D vssd1 vssd1 vccd1 vccd1 _5305_/X sky130_fd_sc_hd__and4_1
XFILLER_88_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8024_ _8024_/A _8098_/A vssd1 vssd1 vccd1 vccd1 _8028_/A sky130_fd_sc_hd__nand2_2
X_5236_ _4950_/X _5228_/X _5235_/Y _5263_/A _5259_/C vssd1 vssd1 vccd1 vccd1 _5236_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_84_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5167_ _4715_/B _5263_/C _4969_/A _5166_/X vssd1 vssd1 vccd1 vccd1 _5168_/B sky130_fd_sc_hd__o31a_1
XFILLER_96_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5098_ _5135_/A _5098_/B _5098_/C _5135_/C vssd1 vssd1 vccd1 vccd1 _5098_/X sky130_fd_sc_hd__or4_1
X_8926_ _8926_/A _4412_/Y vssd1 vssd1 vccd1 vccd1 io_out[13] sky130_fd_sc_hd__ebufn_8
XFILLER_83_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7808_ _7794_/A _8660_/Q _7799_/A _7799_/B _7722_/A vssd1 vssd1 vccd1 vccd1 _7809_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_52_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7739_ _7739_/A _7739_/B vssd1 vssd1 vccd1 vccd1 _7821_/B sky130_fd_sc_hd__nand2_1
XFILLER_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6070_ _6070_/A _6264_/A vssd1 vssd1 vccd1 vccd1 _6093_/B sky130_fd_sc_hd__nor2_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5021_ _5172_/C vssd1 vssd1 vccd1 vccd1 _5250_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_38_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8711_ _8720_/CLK _8711_/D vssd1 vssd1 vccd1 vccd1 _8711_/Q sky130_fd_sc_hd__dfxtp_1
X_6972_ _7079_/A _7079_/B _6980_/B _6971_/B _6971_/A vssd1 vssd1 vccd1 vccd1 _7090_/A
+ sky130_fd_sc_hd__a32o_1
X_5923_ _5922_/A _6144_/A _5922_/D _5922_/C vssd1 vssd1 vccd1 vccd1 _5923_/X sky130_fd_sc_hd__a31o_1
X_5854_ _5773_/A _5775_/A _5920_/A vssd1 vssd1 vccd1 vccd1 _5932_/A sky130_fd_sc_hd__mux2_2
X_8642_ _8723_/CLK _8642_/D vssd1 vssd1 vccd1 vccd1 _8642_/Q sky130_fd_sc_hd__dfxtp_1
X_8573_ _8578_/B _8573_/B _7887_/Y vssd1 vssd1 vccd1 vccd1 _8573_/X sky130_fd_sc_hd__or3b_2
XFILLER_21_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4805_ _7642_/A _4805_/B _4809_/B vssd1 vssd1 vccd1 vccd1 _4806_/A sky130_fd_sc_hd__and3_1
X_5785_ _5851_/C _5785_/B vssd1 vssd1 vccd1 vccd1 _5786_/B sky130_fd_sc_hd__xnor2_1
X_7524_ _7522_/X _7523_/Y _7524_/S vssd1 vssd1 vccd1 vccd1 _7540_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4736_ _4736_/A vssd1 vssd1 vccd1 vccd1 _5130_/A sky130_fd_sc_hd__clkbuf_2
X_4667_ _4670_/C _4667_/B vssd1 vssd1 vccd1 vccd1 _8646_/D sky130_fd_sc_hd__nor2_1
X_7455_ _7455_/A _7455_/B vssd1 vssd1 vccd1 vccd1 _7456_/B sky130_fd_sc_hd__xnor2_1
X_6406_ _6406_/A _6406_/B vssd1 vssd1 vccd1 vccd1 _6407_/B sky130_fd_sc_hd__nand2_1
X_7386_ _7378_/A _7309_/B _7305_/B _7385_/X vssd1 vssd1 vccd1 vccd1 _7387_/B sky130_fd_sc_hd__a31oi_2
X_6337_ _6337_/A _6337_/B vssd1 vssd1 vccd1 vccd1 _6338_/B sky130_fd_sc_hd__xnor2_1
X_4598_ _4598_/A vssd1 vssd1 vccd1 vccd1 _8932_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_1_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6268_ _6268_/A _6268_/B _6268_/C vssd1 vssd1 vccd1 vccd1 _6269_/B sky130_fd_sc_hd__or3_1
X_8007_ _8157_/A vssd1 vssd1 vccd1 vccd1 _8371_/A sky130_fd_sc_hd__clkbuf_2
X_6199_ _6260_/B _6199_/B vssd1 vssd1 vccd1 vccd1 _6205_/A sky130_fd_sc_hd__xnor2_1
XFILLER_69_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5219_ _5219_/A _5219_/B vssd1 vssd1 vccd1 vccd1 _5219_/X sky130_fd_sc_hd__or2_1
XFILLER_28_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8909_ _8909_/A _4392_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[28] sky130_fd_sc_hd__ebufn_8
XFILLER_44_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5570_ _8721_/Q _8658_/Q vssd1 vssd1 vccd1 vccd1 _5572_/A sky130_fd_sc_hd__and2b_1
X_4521_ _6627_/B vssd1 vssd1 vccd1 vccd1 _7679_/A sky130_fd_sc_hd__buf_2
X_4452_ _4456_/A vssd1 vssd1 vccd1 vccd1 _4452_/Y sky130_fd_sc_hd__inv_2
X_7240_ _7240_/A _7240_/B vssd1 vssd1 vccd1 vccd1 _7253_/A sky130_fd_sc_hd__xnor2_1
XFILLER_104_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4383_ _4395_/A vssd1 vssd1 vccd1 vccd1 _4388_/A sky130_fd_sc_hd__clkbuf_2
X_7171_ _6966_/B _7417_/A _7400_/A vssd1 vssd1 vccd1 vccd1 _7179_/A sky130_fd_sc_hd__a21oi_1
X_6122_ _6122_/A _6122_/B vssd1 vssd1 vccd1 vccd1 _6123_/B sky130_fd_sc_hd__xnor2_2
XFILLER_98_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6053_ _6053_/A _6030_/B vssd1 vssd1 vccd1 vccd1 _6053_/X sky130_fd_sc_hd__or2b_1
XFILLER_85_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5004_ _5004_/A vssd1 vssd1 vccd1 vccd1 _5159_/B sky130_fd_sc_hd__clkbuf_2
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6955_ _6955_/A _6992_/B vssd1 vssd1 vccd1 vccd1 _6956_/B sky130_fd_sc_hd__xnor2_1
XFILLER_81_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5906_ _5973_/B _5906_/B vssd1 vssd1 vccd1 vccd1 _5911_/A sky130_fd_sc_hd__xnor2_2
XFILLER_22_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8625_ _8784_/Q _7644_/X _8624_/Y vssd1 vssd1 vccd1 vccd1 _8784_/D sky130_fd_sc_hd__a21o_1
X_6886_ _6886_/A _6886_/B vssd1 vssd1 vccd1 vccd1 _6887_/B sky130_fd_sc_hd__xor2_1
XFILLER_34_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5837_ _5837_/A _5837_/B vssd1 vssd1 vccd1 vccd1 _5838_/B sky130_fd_sc_hd__xnor2_1
X_5768_ _5852_/A _5913_/A vssd1 vssd1 vccd1 vccd1 _5783_/A sky130_fd_sc_hd__nand2_1
X_8556_ _8556_/A _8556_/B vssd1 vssd1 vccd1 vccd1 _8558_/A sky130_fd_sc_hd__xnor2_1
XFILLER_22_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8487_ _8487_/A _8487_/B vssd1 vssd1 vccd1 vccd1 _8490_/A sky130_fd_sc_hd__xnor2_1
X_4719_ _4719_/A vssd1 vssd1 vccd1 vccd1 _8653_/D sky130_fd_sc_hd__clkbuf_1
X_7507_ _7508_/A _7508_/B vssd1 vssd1 vccd1 vccd1 _7507_/Y sky130_fd_sc_hd__nand2_1
X_5699_ _6147_/A _5853_/A vssd1 vssd1 vccd1 vccd1 _5700_/C sky130_fd_sc_hd__nand2_1
X_7438_ _7438_/A _7438_/B vssd1 vssd1 vccd1 vccd1 _7438_/X sky130_fd_sc_hd__and2_1
X_7369_ _7462_/A _7462_/B vssd1 vssd1 vccd1 vccd1 _7482_/B sky130_fd_sc_hd__xor2_1
XFILLER_89_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6740_ _6732_/X _6775_/B _6755_/B vssd1 vssd1 vccd1 vccd1 _6770_/A sky130_fd_sc_hd__a21oi_4
XFILLER_90_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6671_ _7030_/A _6671_/B vssd1 vssd1 vccd1 vccd1 _6725_/B sky130_fd_sc_hd__or2_1
X_8410_ _8345_/A _8345_/B _8409_/X vssd1 vssd1 vccd1 vccd1 _8475_/A sky130_fd_sc_hd__a21oi_1
X_5622_ _5608_/A _5608_/B _5615_/X vssd1 vssd1 vccd1 vccd1 _5634_/C sky130_fd_sc_hd__a21o_1
X_8341_ _8341_/A _8341_/B vssd1 vssd1 vccd1 vccd1 _8342_/B sky130_fd_sc_hd__nand2_1
X_5553_ _5700_/A vssd1 vssd1 vccd1 vccd1 _5766_/A sky130_fd_sc_hd__clkbuf_2
X_4504_ _6653_/B vssd1 vssd1 vccd1 vccd1 _6673_/B sky130_fd_sc_hd__clkbuf_4
X_8272_ _8272_/A _8272_/B _8272_/C _8272_/D vssd1 vssd1 vccd1 vccd1 _8279_/B sky130_fd_sc_hd__or4_1
X_5484_ _5484_/A _5484_/B vssd1 vssd1 vccd1 vccd1 _5484_/X sky130_fd_sc_hd__or2_1
X_4435_ _4438_/A vssd1 vssd1 vccd1 vccd1 _4435_/Y sky130_fd_sc_hd__inv_2
X_7223_ _7223_/A _7042_/B vssd1 vssd1 vccd1 vccd1 _7223_/X sky130_fd_sc_hd__or2b_1
X_4366_ _4369_/A vssd1 vssd1 vccd1 vccd1 _4366_/Y sky130_fd_sc_hd__inv_2
X_7154_ _7133_/B _7154_/B vssd1 vssd1 vccd1 vccd1 _7154_/X sky130_fd_sc_hd__and2b_1
X_6105_ _6137_/A _6137_/B vssd1 vssd1 vccd1 vccd1 _6123_/A sky130_fd_sc_hd__xor2_2
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7085_ _7086_/B _7086_/A vssd1 vssd1 vccd1 vccd1 _7092_/A sky130_fd_sc_hd__or2b_1
X_6036_ _6036_/A _6036_/B _6036_/C vssd1 vssd1 vccd1 vccd1 _6036_/Y sky130_fd_sc_hd__nor3_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7987_ _8006_/B vssd1 vssd1 vccd1 vccd1 _8172_/B sky130_fd_sc_hd__clkbuf_2
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6938_ _6938_/A _6938_/B vssd1 vssd1 vccd1 vccd1 _6939_/B sky130_fd_sc_hd__xnor2_1
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6869_ _6883_/A _6869_/B _6869_/C vssd1 vssd1 vccd1 vccd1 _6871_/A sky130_fd_sc_hd__and3_1
X_8608_ _8608_/A _8614_/B vssd1 vssd1 vccd1 vccd1 _8609_/B sky130_fd_sc_hd__xnor2_1
XFILLER_10_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8539_ _8539_/A _8539_/B vssd1 vssd1 vccd1 vccd1 _8539_/Y sky130_fd_sc_hd__nand2_1
XFILLER_10_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7910_ _7910_/A _7910_/B _7910_/C vssd1 vssd1 vccd1 vccd1 _7919_/A sky130_fd_sc_hd__nand3_1
X_8890_ _8890_/A _4368_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[9] sky130_fd_sc_hd__ebufn_8
XFILLER_48_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7841_ _8774_/Q _7842_/B vssd1 vssd1 vccd1 vccd1 _8102_/A sky130_fd_sc_hd__or2_1
XFILLER_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7772_ _7772_/A _7772_/B vssd1 vssd1 vccd1 vccd1 _7773_/C sky130_fd_sc_hd__and2_1
X_4984_ _5215_/B _5228_/A _5142_/C vssd1 vssd1 vccd1 vccd1 _5199_/A sky130_fd_sc_hd__nor3_2
X_6723_ _6958_/A _7078_/B _6959_/B vssd1 vssd1 vccd1 vccd1 _6723_/X sky130_fd_sc_hd__and3_1
X_6654_ _7794_/B _7583_/A vssd1 vssd1 vccd1 vccd1 _6678_/A sky130_fd_sc_hd__or2b_2
X_5605_ _5732_/A _5732_/B vssd1 vssd1 vccd1 vccd1 _5727_/B sky130_fd_sc_hd__xor2_1
XFILLER_31_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6585_ _6580_/A _6580_/B _6578_/B vssd1 vssd1 vccd1 vccd1 _6586_/B sky130_fd_sc_hd__a21oi_1
X_8324_ _8568_/B _8289_/B _8292_/B _8323_/Y vssd1 vssd1 vccd1 vccd1 _8425_/B sky130_fd_sc_hd__a31o_1
X_5536_ _5683_/A _5683_/B vssd1 vssd1 vccd1 vccd1 _5684_/A sky130_fd_sc_hd__nor2_1
X_8255_ _8362_/A _8255_/B vssd1 vssd1 vccd1 vccd1 _8284_/A sky130_fd_sc_hd__and2_1
X_5467_ _5467_/A _5467_/B vssd1 vssd1 vccd1 vccd1 _5467_/Y sky130_fd_sc_hd__nor2_1
X_4418_ _4419_/A vssd1 vssd1 vccd1 vccd1 _4418_/Y sky130_fd_sc_hd__inv_2
X_7206_ _7380_/A _7300_/A vssd1 vssd1 vccd1 vccd1 _7306_/B sky130_fd_sc_hd__xnor2_1
X_8186_ _8244_/A _8186_/B vssd1 vssd1 vccd1 vccd1 _8187_/B sky130_fd_sc_hd__nor2_2
X_5398_ _8699_/Q _5401_/C vssd1 vssd1 vccd1 vccd1 _5400_/A sky130_fd_sc_hd__and2_1
XFILLER_98_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7137_ _7137_/A _7137_/B vssd1 vssd1 vccd1 vccd1 _7151_/B sky130_fd_sc_hd__xor2_1
XFILLER_59_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7068_ _7068_/A _7068_/B vssd1 vssd1 vccd1 vccd1 _7525_/A sky130_fd_sc_hd__nor2_1
X_6019_ _6019_/A _6019_/B vssd1 vssd1 vccd1 vccd1 _6057_/A sky130_fd_sc_hd__xor2_1
XFILLER_46_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6370_ _6370_/A _6370_/B vssd1 vssd1 vccd1 vccd1 _6372_/A sky130_fd_sc_hd__xnor2_1
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5321_ _8677_/Q _5326_/B vssd1 vssd1 vccd1 vccd1 _5321_/X sky130_fd_sc_hd__or2_1
X_8040_ _8058_/A _8039_/B _8039_/C vssd1 vssd1 vccd1 vccd1 _8040_/Y sky130_fd_sc_hd__o21ai_1
X_5252_ _5197_/D _5154_/X _5156_/X _4702_/D _5251_/X vssd1 vssd1 vccd1 vccd1 _5252_/X
+ sky130_fd_sc_hd__o221a_1
X_5183_ _5183_/A vssd1 vssd1 vccd1 vccd1 _5274_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_68_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8942_ _8942_/A _4431_/Y vssd1 vssd1 vccd1 vccd1 io_out[29] sky130_fd_sc_hd__ebufn_8
XFILLER_49_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7824_ _8262_/A vssd1 vssd1 vccd1 vccd1 _8382_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7755_ _8450_/B _8182_/A _7768_/A vssd1 vssd1 vccd1 vccd1 _7755_/X sky130_fd_sc_hd__or3b_2
XFILLER_51_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4967_ _5148_/A _5234_/A vssd1 vssd1 vccd1 vccd1 _4967_/X sky130_fd_sc_hd__or2_1
X_7686_ _7684_/X _7686_/B vssd1 vssd1 vccd1 vccd1 _7688_/C sky130_fd_sc_hd__and2b_1
X_6706_ _7392_/A vssd1 vssd1 vccd1 vccd1 _7120_/B sky130_fd_sc_hd__clkbuf_2
X_4898_ _4910_/A _4925_/A vssd1 vssd1 vccd1 vccd1 _5074_/B sky130_fd_sc_hd__nor2_1
X_6637_ _6648_/A _6637_/B vssd1 vssd1 vccd1 vccd1 _6671_/B sky130_fd_sc_hd__xnor2_1
X_6568_ _6568_/A vssd1 vssd1 vccd1 vccd1 _6569_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_98_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8307_ _8317_/A _8317_/B vssd1 vssd1 vccd1 vccd1 _8308_/B sky130_fd_sc_hd__xor2_2
X_5519_ _7700_/A _8711_/Q vssd1 vssd1 vccd1 vccd1 _5544_/A sky130_fd_sc_hd__or2b_1
XFILLER_3_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6499_ _6501_/B _6499_/B _6517_/B vssd1 vssd1 vccd1 vccd1 _6500_/A sky130_fd_sc_hd__and3b_1
X_8238_ _8238_/A vssd1 vssd1 vccd1 vccd1 _8527_/A sky130_fd_sc_hd__clkbuf_2
X_8169_ _8169_/A _8169_/B vssd1 vssd1 vccd1 vccd1 _8256_/B sky130_fd_sc_hd__xnor2_2
XFILLER_78_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5870_ _5867_/X _5868_/Y _5810_/X _5792_/X vssd1 vssd1 vccd1 vccd1 _5875_/B sky130_fd_sc_hd__a211o_1
X_4821_ _8664_/Q _8663_/Q _7672_/B vssd1 vssd1 vccd1 vccd1 _4850_/C sky130_fd_sc_hd__o21a_1
XFILLER_33_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4752_ _4760_/A _4752_/B _4758_/C vssd1 vssd1 vccd1 vccd1 _4753_/A sky130_fd_sc_hd__and3_1
XFILLER_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7540_ _7540_/A _7540_/B _7540_/C _7539_/X vssd1 vssd1 vccd1 vccd1 _7540_/X sky130_fd_sc_hd__or4b_1
X_4683_ _5462_/A _4679_/C _5440_/C vssd1 vssd1 vccd1 vccd1 _4684_/B sky130_fd_sc_hd__o21ai_1
X_7471_ _7471_/A _7471_/B vssd1 vssd1 vccd1 vccd1 _7472_/B sky130_fd_sc_hd__xnor2_1
X_6422_ _6423_/A _6423_/B _6423_/C _6423_/D vssd1 vssd1 vccd1 vccd1 _6422_/Y sky130_fd_sc_hd__o22ai_1
X_6353_ _6353_/A _6353_/B vssd1 vssd1 vccd1 vccd1 _6354_/B sky130_fd_sc_hd__xnor2_1
X_6284_ _6284_/A _6284_/B vssd1 vssd1 vccd1 vccd1 _6300_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5304_ _4543_/A _4568_/B _5302_/Y _5303_/X vssd1 vssd1 vccd1 vccd1 _5305_/D sky130_fd_sc_hd__o211a_1
X_8023_ _7955_/A _8023_/B vssd1 vssd1 vccd1 vccd1 _8030_/B sky130_fd_sc_hd__and2b_1
X_5235_ _5235_/A vssd1 vssd1 vccd1 vccd1 _5235_/Y sky130_fd_sc_hd__inv_2
X_5166_ _5188_/A _5192_/B _5190_/A _5118_/B vssd1 vssd1 vccd1 vccd1 _5166_/X sky130_fd_sc_hd__or4b_1
XFILLER_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5097_ _5154_/A _5119_/A vssd1 vssd1 vccd1 vccd1 _5135_/C sky130_fd_sc_hd__or2_1
X_8925_ _8925_/A _4411_/Y vssd1 vssd1 vccd1 vccd1 io_out[12] sky130_fd_sc_hd__ebufn_8
XFILLER_17_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5999_ _6075_/B _5999_/B vssd1 vssd1 vccd1 vccd1 _6000_/B sky130_fd_sc_hd__nor2_1
X_7807_ _8381_/A _7807_/B vssd1 vssd1 vccd1 vccd1 _7813_/B sky130_fd_sc_hd__and2b_1
XFILLER_52_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7738_ _8595_/A vssd1 vssd1 vccd1 vccd1 _7739_/A sky130_fd_sc_hd__inv_2
X_7669_ _7943_/A _7667_/Y _7668_/Y vssd1 vssd1 vccd1 vccd1 _8774_/D sky130_fd_sc_hd__a21oi_1
XFILLER_3_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5020_ _5042_/A _5209_/B vssd1 vssd1 vccd1 vccd1 _5031_/B sky130_fd_sc_hd__or2_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6971_ _6971_/A _6971_/B vssd1 vssd1 vccd1 vccd1 _6980_/B sky130_fd_sc_hd__xor2_1
X_8710_ _8765_/CLK _8710_/D vssd1 vssd1 vccd1 vccd1 _8710_/Q sky130_fd_sc_hd__dfxtp_1
X_5922_ _5922_/A _6144_/A _5922_/C _5922_/D vssd1 vssd1 vccd1 vccd1 _6036_/A sky130_fd_sc_hd__and4_1
X_5853_ _5853_/A _5853_/B vssd1 vssd1 vccd1 vccd1 _5920_/A sky130_fd_sc_hd__or2_2
XFILLER_61_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8641_ _8723_/CLK _8641_/D vssd1 vssd1 vccd1 vccd1 _8641_/Q sky130_fd_sc_hd__dfxtp_1
X_5784_ _5872_/B _5784_/B vssd1 vssd1 vccd1 vccd1 _5785_/B sky130_fd_sc_hd__nor2_1
X_8572_ _7888_/A _8577_/B _7979_/X vssd1 vssd1 vccd1 vccd1 _8573_/B sky130_fd_sc_hd__a21bo_1
XFILLER_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4804_ _4804_/A _4804_/B _4804_/C vssd1 vssd1 vccd1 vccd1 _4809_/B sky130_fd_sc_hd__nand3_1
X_4735_ _4973_/A _4973_/B vssd1 vssd1 vccd1 vccd1 _4736_/A sky130_fd_sc_hd__nor2_1
XFILLER_9_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7523_ _7523_/A _7523_/B vssd1 vssd1 vccd1 vccd1 _7523_/Y sky130_fd_sc_hd__nand2_1
X_4666_ _8646_/Q _4665_/B _4640_/X vssd1 vssd1 vccd1 vccd1 _4667_/B sky130_fd_sc_hd__o21ai_1
X_7454_ _7454_/A _7454_/B vssd1 vssd1 vccd1 vccd1 _7455_/B sky130_fd_sc_hd__xnor2_1
X_6405_ _6405_/A _8705_/Q vssd1 vssd1 vccd1 vccd1 _6406_/B sky130_fd_sc_hd__or2b_1
X_4597_ _8678_/Q _5305_/A vssd1 vssd1 vccd1 vccd1 _4598_/A sky130_fd_sc_hd__and2_1
X_7385_ _7304_/B _7485_/B vssd1 vssd1 vccd1 vccd1 _7385_/X sky130_fd_sc_hd__and2b_1
X_6336_ _6336_/A _6336_/B vssd1 vssd1 vccd1 vccd1 _6337_/B sky130_fd_sc_hd__xnor2_1
XFILLER_88_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6267_ _6268_/A _6268_/B _6268_/C vssd1 vssd1 vccd1 vccd1 _6269_/A sky130_fd_sc_hd__o21ai_1
X_8006_ _8568_/C _8006_/B vssd1 vssd1 vccd1 vccd1 _8157_/A sky130_fd_sc_hd__nor2_2
XFILLER_76_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6198_ _5994_/B _6275_/S _6197_/Y _6085_/A vssd1 vssd1 vccd1 vccd1 _6199_/B sky130_fd_sc_hd__o2bb2a_1
X_5218_ _4715_/B _5221_/B _5174_/A _5188_/D _5215_/X vssd1 vssd1 vccd1 vccd1 _5219_/B
+ sky130_fd_sc_hd__o32a_1
XFILLER_56_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5149_ _5250_/C _5149_/B _5149_/C _5149_/D vssd1 vssd1 vccd1 vccd1 _5150_/B sky130_fd_sc_hd__nor4_1
XFILLER_84_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8908_ _8908_/A _4391_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[27] sky130_fd_sc_hd__ebufn_8
XFILLER_71_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4520_ _8667_/Q vssd1 vssd1 vccd1 vccd1 _6627_/B sky130_fd_sc_hd__clkbuf_2
X_4451_ _4457_/A vssd1 vssd1 vccd1 vccd1 _4456_/A sky130_fd_sc_hd__buf_6
X_7170_ _7024_/A _7024_/B _7169_/X vssd1 vssd1 vccd1 vccd1 _7259_/A sky130_fd_sc_hd__o21a_1
X_6121_ _6121_/A _6121_/B vssd1 vssd1 vccd1 vccd1 _6122_/B sky130_fd_sc_hd__nand2_1
XFILLER_98_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4382_ _4382_/A vssd1 vssd1 vccd1 vccd1 _4382_/Y sky130_fd_sc_hd__inv_2
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6052_ _6044_/A _6044_/B _6043_/A vssd1 vssd1 vccd1 vccd1 _6125_/A sky130_fd_sc_hd__o21ai_2
XFILLER_98_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5003_ _5172_/A vssd1 vssd1 vccd1 vccd1 _5215_/A sky130_fd_sc_hd__clkbuf_2
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6954_ _6954_/A _6954_/B vssd1 vssd1 vccd1 vccd1 _6992_/B sky130_fd_sc_hd__xor2_1
X_5905_ _5905_/A _5905_/B vssd1 vssd1 vccd1 vccd1 _5906_/B sky130_fd_sc_hd__xnor2_1
X_8624_ _7644_/X _8623_/Y _7624_/X vssd1 vssd1 vccd1 vccd1 _8624_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_14_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6885_ _6885_/A _6885_/B vssd1 vssd1 vccd1 vccd1 _6886_/B sky130_fd_sc_hd__xnor2_1
XFILLER_22_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5836_ _5741_/A _5751_/A _5743_/B _5743_/A vssd1 vssd1 vccd1 vccd1 _5907_/A sky130_fd_sc_hd__a22o_1
X_5767_ _5662_/B _5657_/B _5766_/X vssd1 vssd1 vccd1 vccd1 _5779_/A sky130_fd_sc_hd__a21oi_1
X_8555_ _8554_/B _8563_/A _8554_/A vssd1 vssd1 vccd1 vccd1 _8555_/Y sky130_fd_sc_hd__o21ai_1
X_5698_ _5698_/A _6107_/A vssd1 vssd1 vccd1 vccd1 _5926_/A sky130_fd_sc_hd__nand2_1
X_8486_ _8479_/A _8484_/B _8479_/B vssd1 vssd1 vccd1 vccd1 _8547_/B sky130_fd_sc_hd__a21bo_1
X_4718_ _4760_/A _4718_/B _4745_/A vssd1 vssd1 vccd1 vccd1 _4719_/A sky130_fd_sc_hd__and3_1
X_7506_ _7430_/A _7430_/B _7505_/X vssd1 vssd1 vccd1 vccd1 _7510_/A sky130_fd_sc_hd__a21oi_1
X_7437_ _7438_/A _7438_/B vssd1 vssd1 vccd1 vccd1 _7437_/X sky130_fd_sc_hd__or2_1
XFILLER_30_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4649_ _4652_/C _4649_/B vssd1 vssd1 vccd1 vccd1 _8640_/D sky130_fd_sc_hd__nor2_1
X_8875__92 vssd1 vssd1 vccd1 vccd1 _8875__92/HI _8984_/A sky130_fd_sc_hd__conb_1
XFILLER_89_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7368_ _7461_/A _7461_/B vssd1 vssd1 vccd1 vccd1 _7462_/B sky130_fd_sc_hd__xor2_1
XFILLER_103_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6319_ _6279_/A _6280_/A _6279_/B vssd1 vssd1 vccd1 vccd1 _6320_/B sky130_fd_sc_hd__o21ba_1
X_7299_ _6966_/B _7176_/B _7405_/A _7412_/A vssd1 vssd1 vccd1 vccd1 _7318_/A sky130_fd_sc_hd__o211ai_2
XFILLER_39_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6670_ _6670_/A _6670_/B vssd1 vssd1 vccd1 vccd1 _7030_/A sky130_fd_sc_hd__xnor2_4
X_5621_ _7794_/B _6427_/A vssd1 vssd1 vccd1 vccd1 _5634_/A sky130_fd_sc_hd__or2b_2
XFILLER_31_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8340_ _8340_/A _8296_/B vssd1 vssd1 vccd1 vccd1 _8341_/B sky130_fd_sc_hd__or2b_1
X_5552_ _5552_/A _5552_/B vssd1 vssd1 vccd1 vccd1 _5700_/A sky130_fd_sc_hd__nand2_1
X_8271_ _8463_/A vssd1 vssd1 vccd1 vccd1 _8279_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4503_ _8661_/Q vssd1 vssd1 vccd1 vccd1 _6653_/B sky130_fd_sc_hd__buf_2
XFILLER_8_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5483_ _8713_/Q vssd1 vssd1 vccd1 vccd1 _5648_/A sky130_fd_sc_hd__inv_2
X_4434_ _4438_/A vssd1 vssd1 vccd1 vccd1 _4434_/Y sky130_fd_sc_hd__inv_2
X_7222_ _7373_/A _7058_/B _7221_/Y vssd1 vssd1 vccd1 vccd1 _7256_/A sky130_fd_sc_hd__o21a_1
X_4365_ _4369_/A vssd1 vssd1 vccd1 vccd1 _4365_/Y sky130_fd_sc_hd__inv_2
X_7153_ _7151_/A _7151_/B _7516_/A vssd1 vssd1 vccd1 vccd1 _7519_/B sky130_fd_sc_hd__a21o_1
X_6104_ _6104_/A _6104_/B vssd1 vssd1 vccd1 vccd1 _6137_/B sky130_fd_sc_hd__xnor2_2
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7084_ _7098_/A _7098_/B _7083_/Y vssd1 vssd1 vccd1 vccd1 _7086_/A sky130_fd_sc_hd__a21bo_1
X_6035_ _6249_/A _6059_/A vssd1 vssd1 vccd1 vccd1 _6036_/C sky130_fd_sc_hd__nor2_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7986_ _8008_/A _7908_/B _7908_/C vssd1 vssd1 vccd1 vccd1 _7994_/A sky130_fd_sc_hd__a21bo_1
XFILLER_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6937_ _7228_/B _6937_/B vssd1 vssd1 vccd1 vccd1 _6938_/B sky130_fd_sc_hd__xor2_1
XFILLER_25_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6868_ _6873_/A _6873_/B _7176_/A vssd1 vssd1 vccd1 vccd1 _6869_/C sky130_fd_sc_hd__o21ai_1
X_5819_ _5892_/A _6192_/A _5819_/C _5819_/D vssd1 vssd1 vccd1 vccd1 _5890_/A sky130_fd_sc_hd__or4_1
X_8607_ _8602_/A _8602_/B _8600_/A vssd1 vssd1 vccd1 vccd1 _8614_/B sky130_fd_sc_hd__a21oi_1
XFILLER_10_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8538_ _8538_/A _8538_/B vssd1 vssd1 vccd1 vccd1 _8543_/A sky130_fd_sc_hd__xnor2_1
XFILLER_10_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6799_ _6799_/A _7303_/A vssd1 vssd1 vccd1 vccd1 _6801_/C sky130_fd_sc_hd__xnor2_1
XFILLER_22_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8469_ _8469_/A _8469_/B vssd1 vssd1 vccd1 vccd1 _8470_/B sky130_fd_sc_hd__nor2_1
XFILLER_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7840_ _7784_/A _7784_/B _7839_/X vssd1 vssd1 vccd1 vccd1 _7938_/A sky130_fd_sc_hd__a21oi_2
XFILLER_36_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7771_ _7772_/A _7772_/B vssd1 vssd1 vccd1 vccd1 _7872_/B sky130_fd_sc_hd__nor2_1
XFILLER_51_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4983_ _5153_/C vssd1 vssd1 vccd1 vccd1 _5228_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_23_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6722_ _6729_/A _6722_/B vssd1 vssd1 vccd1 vccd1 _6959_/B sky130_fd_sc_hd__and2_1
XFILLER_23_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6653_ _6653_/A _6653_/B vssd1 vssd1 vccd1 vccd1 _6674_/B sky130_fd_sc_hd__or2_1
XFILLER_31_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5604_ _5608_/A _5608_/B _5615_/A vssd1 vssd1 vccd1 vccd1 _5732_/B sky130_fd_sc_hd__a21oi_2
X_6584_ _6582_/Y _6584_/B vssd1 vssd1 vccd1 vccd1 _6586_/A sky130_fd_sc_hd__and2b_1
X_8323_ _8487_/A _8323_/B vssd1 vssd1 vccd1 vccd1 _8323_/Y sky130_fd_sc_hd__nor2_1
X_5535_ _5681_/A _5535_/B vssd1 vssd1 vccd1 vccd1 _5683_/B sky130_fd_sc_hd__xnor2_1
XFILLER_11_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8254_ _8254_/A _8254_/B _8254_/C vssd1 vssd1 vccd1 vccd1 _8255_/B sky130_fd_sc_hd__or3_1
X_5466_ _5458_/B _5460_/B _5458_/A vssd1 vssd1 vccd1 vccd1 _5467_/B sky130_fd_sc_hd__o21ba_1
X_4417_ _4419_/A vssd1 vssd1 vccd1 vccd1 _4417_/Y sky130_fd_sc_hd__inv_2
X_7205_ _7302_/A _7205_/B vssd1 vssd1 vccd1 vccd1 _7300_/A sky130_fd_sc_hd__nor2_2
X_8185_ _8185_/A _8185_/B _8453_/A vssd1 vssd1 vccd1 vccd1 _8186_/B sky130_fd_sc_hd__and3_1
X_8845__62 vssd1 vssd1 vccd1 vccd1 _8845__62/HI _8954_/A sky130_fd_sc_hd__conb_1
XFILLER_59_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5397_ _5401_/C _5397_/B vssd1 vssd1 vccd1 vccd1 _8698_/D sky130_fd_sc_hd__nor2_1
X_7136_ _7138_/A _7138_/B vssd1 vssd1 vccd1 vccd1 _7151_/A sky130_fd_sc_hd__and2_1
X_7067_ _7067_/A _7067_/B _7067_/C vssd1 vssd1 vccd1 vccd1 _7068_/B sky130_fd_sc_hd__and3_1
X_6018_ _5861_/B _6251_/A _6171_/A _6017_/Y vssd1 vssd1 vccd1 vccd1 _6019_/B sky130_fd_sc_hd__a31o_1
XFILLER_86_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7969_ _7970_/A _7970_/B vssd1 vssd1 vccd1 vccd1 _8051_/A sky130_fd_sc_hd__or2_1
XFILLER_27_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5320_ _5320_/A vssd1 vssd1 vccd1 vccd1 _5320_/X sky130_fd_sc_hd__clkbuf_2
X_5251_ _5251_/A _5251_/B _5251_/C vssd1 vssd1 vccd1 vccd1 _5251_/X sky130_fd_sc_hd__or3_1
XFILLER_87_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5182_ _5182_/A _5266_/B vssd1 vssd1 vccd1 vccd1 _5291_/C sky130_fd_sc_hd__nand2_2
XFILLER_95_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8941_ _8941_/A _4430_/Y vssd1 vssd1 vccd1 vccd1 io_out[28] sky130_fd_sc_hd__ebufn_8
XFILLER_95_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7823_ _7826_/A _7902_/B _7828_/B vssd1 vssd1 vccd1 vccd1 _8262_/A sky130_fd_sc_hd__and3_1
XFILLER_51_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7754_ _7754_/A _8172_/A vssd1 vssd1 vccd1 vccd1 _7768_/A sky130_fd_sc_hd__nand2_1
X_6705_ _7034_/B vssd1 vssd1 vccd1 vccd1 _7392_/A sky130_fd_sc_hd__clkbuf_2
X_4966_ _4966_/A vssd1 vssd1 vccd1 vccd1 _5234_/A sky130_fd_sc_hd__clkbuf_2
X_7685_ _7685_/A _8771_/Q vssd1 vssd1 vccd1 vccd1 _7686_/B sky130_fd_sc_hd__or2b_1
XFILLER_22_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4897_ _4901_/A _4897_/B _4897_/C _4778_/A vssd1 vssd1 vccd1 vccd1 _4925_/A sky130_fd_sc_hd__or4b_4
X_6636_ _6898_/A _6774_/A vssd1 vssd1 vccd1 vccd1 _7186_/B sky130_fd_sc_hd__nand2_1
X_6567_ _6567_/A vssd1 vssd1 vccd1 vccd1 _6567_/X sky130_fd_sc_hd__clkbuf_2
X_8306_ _8306_/A _8306_/B vssd1 vssd1 vccd1 vccd1 _8317_/B sky130_fd_sc_hd__xnor2_2
X_5518_ _8711_/Q _8669_/Q vssd1 vssd1 vccd1 vccd1 _5518_/X sky130_fd_sc_hd__and2b_1
Xclkbuf_4_1_0_wb_clk_i clkbuf_4_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _8732_/CLK
+ sky130_fd_sc_hd__clkbuf_2
X_6498_ _6497_/B _8734_/Q _6491_/A _8736_/Q vssd1 vssd1 vccd1 vccd1 _6499_/B sky130_fd_sc_hd__a31o_1
X_8237_ _8237_/A _8441_/A vssd1 vssd1 vccd1 vccd1 _8245_/A sky130_fd_sc_hd__nand2_1
X_5449_ _5449_/A vssd1 vssd1 vccd1 vccd1 _5449_/X sky130_fd_sc_hd__clkbuf_2
X_8168_ _8272_/C _8272_/D vssd1 vssd1 vccd1 vccd1 _8169_/B sky130_fd_sc_hd__nor2_1
XFILLER_87_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7119_ _7119_/A _7123_/C vssd1 vssd1 vccd1 vccd1 _7119_/X sky130_fd_sc_hd__or2_1
X_8099_ _8099_/A _8327_/A _8099_/C _8099_/D vssd1 vssd1 vccd1 vccd1 _8214_/A sky130_fd_sc_hd__and4_1
XFILLER_86_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4820_ _7672_/B _8664_/Q _8663_/Q _8662_/Q vssd1 vssd1 vccd1 vccd1 _4894_/B sky130_fd_sc_hd__or4b_4
XFILLER_61_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4751_ _5300_/B _4751_/B vssd1 vssd1 vccd1 vccd1 _4758_/C sky130_fd_sc_hd__nand2_1
X_4682_ _5462_/B vssd1 vssd1 vccd1 vccd1 _5440_/C sky130_fd_sc_hd__clkbuf_2
X_7470_ _7470_/A _7470_/B vssd1 vssd1 vccd1 vccd1 _7471_/B sky130_fd_sc_hd__xnor2_1
X_6421_ _6420_/B _6427_/B vssd1 vssd1 vccd1 vccd1 _6423_/D sky130_fd_sc_hd__and2b_1
X_6352_ _6288_/A _6288_/B _6351_/Y vssd1 vssd1 vccd1 vccd1 _6353_/B sky130_fd_sc_hd__o21ai_1
X_6283_ _6346_/A _6283_/B vssd1 vssd1 vccd1 vccd1 _6284_/B sky130_fd_sc_hd__xnor2_1
XFILLER_88_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5303_ _4814_/A _4814_/B _5298_/A _4870_/A _4804_/A vssd1 vssd1 vccd1 vccd1 _5303_/X
+ sky130_fd_sc_hd__o221a_1
X_8815__32 vssd1 vssd1 vccd1 vccd1 _8815__32/HI _8910_/A sky130_fd_sc_hd__conb_1
X_8022_ _7951_/A _8022_/B vssd1 vssd1 vccd1 vccd1 _8113_/A sky130_fd_sc_hd__and2b_1
XFILLER_69_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5234_ _5234_/A _5234_/B vssd1 vssd1 vccd1 vccd1 _5234_/X sky130_fd_sc_hd__or2_1
X_5165_ _5255_/A _5265_/B _4969_/A _5031_/B _5164_/X vssd1 vssd1 vccd1 vccd1 _5165_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_96_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5096_ _5283_/A _5096_/B vssd1 vssd1 vccd1 vccd1 _5098_/C sky130_fd_sc_hd__or2_1
X_8924_ _8924_/A _4410_/Y vssd1 vssd1 vccd1 vccd1 io_out[11] sky130_fd_sc_hd__ebufn_8
XFILLER_17_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7806_ _8661_/Q _7602_/A vssd1 vssd1 vccd1 vccd1 _7807_/B sky130_fd_sc_hd__or2b_2
X_5998_ _6088_/A _5998_/B vssd1 vssd1 vccd1 vccd1 _5999_/B sky130_fd_sc_hd__nor2_1
X_7737_ _7799_/A _7799_/B vssd1 vssd1 vccd1 vccd1 _8155_/A sky130_fd_sc_hd__xor2_4
X_4949_ _5264_/A _5275_/A vssd1 vssd1 vccd1 vccd1 _5251_/B sky130_fd_sc_hd__nand2_1
X_7668_ _7943_/A _7667_/Y _4615_/A vssd1 vssd1 vccd1 vccd1 _7668_/Y sky130_fd_sc_hd__o21ai_1
X_6619_ _7309_/A _7391_/A vssd1 vssd1 vccd1 vccd1 _7120_/A sky130_fd_sc_hd__nand2_2
X_7599_ _7734_/A _8593_/A _8595_/A _7598_/Y vssd1 vssd1 vccd1 vccd1 _7599_/X sky130_fd_sc_hd__a31o_1
XFILLER_3_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6970_ _6970_/A _6970_/B vssd1 vssd1 vccd1 vccd1 _6971_/B sky130_fd_sc_hd__xnor2_1
XFILLER_38_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5921_ _6251_/A _5921_/B vssd1 vssd1 vccd1 vccd1 _5922_/D sky130_fd_sc_hd__or2_1
XFILLER_65_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5852_ _5852_/A _5921_/B vssd1 vssd1 vccd1 vccd1 _5856_/A sky130_fd_sc_hd__nand2_2
XFILLER_80_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8640_ _8730_/CLK _8640_/D vssd1 vssd1 vccd1 vccd1 _8640_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5783_ _5783_/A _5783_/B vssd1 vssd1 vccd1 vccd1 _5784_/B sky130_fd_sc_hd__and2_1
X_8571_ _8571_/A _8571_/B vssd1 vssd1 vccd1 vccd1 _8577_/B sky130_fd_sc_hd__xnor2_1
XFILLER_61_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4803_ _4804_/B _4804_/C _4804_/A vssd1 vssd1 vccd1 vccd1 _4805_/B sky130_fd_sc_hd__a21o_1
X_4734_ _6613_/B _4734_/B vssd1 vssd1 vccd1 vccd1 _4973_/B sky130_fd_sc_hd__nor2_1
X_7522_ _7523_/A _7522_/B vssd1 vssd1 vccd1 vccd1 _7522_/X sky130_fd_sc_hd__or2_1
XFILLER_9_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4665_ _8646_/Q _4665_/B vssd1 vssd1 vccd1 vccd1 _4670_/C sky130_fd_sc_hd__and2_1
X_7453_ _7453_/A _7453_/B vssd1 vssd1 vccd1 vccd1 _7454_/B sky130_fd_sc_hd__xnor2_2
X_4596_ _4596_/A vssd1 vssd1 vccd1 vccd1 _8931_/A sky130_fd_sc_hd__clkbuf_1
X_6404_ _8705_/Q _6405_/A vssd1 vssd1 vccd1 vccd1 _6406_/A sky130_fd_sc_hd__or2b_1
X_7384_ _7384_/A _7384_/B vssd1 vssd1 vccd1 vccd1 _7463_/B sky130_fd_sc_hd__xnor2_2
X_6335_ _6180_/B _6333_/Y _6334_/Y vssd1 vssd1 vccd1 vccd1 _6336_/B sky130_fd_sc_hd__o21a_1
X_8005_ _8061_/B _8004_/C _8004_/A vssd1 vssd1 vccd1 vccd1 _8014_/B sky130_fd_sc_hd__a21o_1
X_6266_ _6323_/A _6266_/B vssd1 vssd1 vccd1 vccd1 _6268_/C sky130_fd_sc_hd__xnor2_1
X_6197_ _6197_/A _6274_/B vssd1 vssd1 vccd1 vccd1 _6197_/Y sky130_fd_sc_hd__nor2_1
XFILLER_57_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5217_ _5176_/A _5163_/B _5214_/X _5216_/X vssd1 vssd1 vccd1 vccd1 _5217_/X sky130_fd_sc_hd__o31a_1
XFILLER_96_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5148_ _5148_/A _5148_/B _5148_/C vssd1 vssd1 vccd1 vccd1 _5148_/X sky130_fd_sc_hd__or3_1
XFILLER_56_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5079_ _5079_/A vssd1 vssd1 vccd1 vccd1 _5261_/D sky130_fd_sc_hd__clkbuf_2
X_8907_ _8907_/A _4390_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[26] sky130_fd_sc_hd__ebufn_8
XFILLER_71_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8769_ _8776_/CLK _8769_/D vssd1 vssd1 vccd1 vccd1 _8769_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_12_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4450_ _4450_/A vssd1 vssd1 vccd1 vccd1 _4450_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4381_ _4382_/A vssd1 vssd1 vccd1 vccd1 _4381_/Y sky130_fd_sc_hd__inv_2
X_6120_ _6120_/A _6120_/B vssd1 vssd1 vccd1 vccd1 _6122_/A sky130_fd_sc_hd__nor2_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6051_ _6047_/A _6047_/B _6050_/Y vssd1 vssd1 vccd1 vccd1 _6293_/A sky130_fd_sc_hd__a21oi_2
XFILLER_98_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5002_ _5077_/B vssd1 vssd1 vccd1 vccd1 _5163_/B sky130_fd_sc_hd__clkbuf_2
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6953_ _6953_/A _6953_/B vssd1 vssd1 vccd1 vccd1 _6954_/B sky130_fd_sc_hd__xnor2_1
XFILLER_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5904_ _6007_/B _5904_/B vssd1 vssd1 vccd1 vccd1 _5905_/B sky130_fd_sc_hd__nand2_1
X_6884_ _6886_/A _7378_/A _6802_/A vssd1 vssd1 vccd1 vccd1 _6885_/B sky130_fd_sc_hd__a21bo_1
XFILLER_34_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5835_ _5835_/A _5897_/A vssd1 vssd1 vccd1 vccd1 _5908_/A sky130_fd_sc_hd__or2_1
X_8623_ _8623_/A _8623_/B vssd1 vssd1 vccd1 vccd1 _8623_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5766_ _5766_/A _5921_/B _5766_/C vssd1 vssd1 vccd1 vccd1 _5766_/X sky130_fd_sc_hd__and3_1
X_8554_ _8554_/A _8554_/B _8563_/A vssd1 vssd1 vccd1 vccd1 _8554_/X sky130_fd_sc_hd__or3_1
XFILLER_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5697_ _5697_/A _5697_/B vssd1 vssd1 vccd1 vccd1 _5710_/A sky130_fd_sc_hd__xnor2_1
X_8485_ _8549_/B _8549_/C _8550_/B _8549_/A vssd1 vssd1 vccd1 vccd1 _8547_/A sky130_fd_sc_hd__a211o_1
X_7505_ _7505_/A _7505_/B vssd1 vssd1 vccd1 vccd1 _7505_/X sky130_fd_sc_hd__and2_1
X_4717_ _4771_/A _5259_/D vssd1 vssd1 vccd1 vccd1 _4745_/A sky130_fd_sc_hd__nand2_1
X_4648_ _8640_/Q _4647_/B _4628_/X vssd1 vssd1 vccd1 vccd1 _4649_/B sky130_fd_sc_hd__o21ai_1
X_7436_ _7438_/A _7438_/B vssd1 vssd1 vccd1 vccd1 _7523_/B sky130_fd_sc_hd__xor2_2
X_4579_ _4579_/A vssd1 vssd1 vccd1 vccd1 _8927_/A sky130_fd_sc_hd__clkbuf_1
X_7367_ _7367_/A _7367_/B vssd1 vssd1 vccd1 vccd1 _7461_/B sky130_fd_sc_hd__xnor2_1
XFILLER_89_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6318_ _6318_/A _6318_/B vssd1 vssd1 vccd1 vccd1 _6341_/A sky130_fd_sc_hd__xnor2_1
X_7298_ _7214_/A _7214_/B _7297_/X vssd1 vssd1 vccd1 vccd1 _7320_/A sky130_fd_sc_hd__a21o_1
XFILLER_103_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6249_ _6249_/A _6252_/B vssd1 vssd1 vccd1 vccd1 _6311_/C sky130_fd_sc_hd__nand2_1
XFILLER_49_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_4_14_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8778_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_82_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5620_ _5620_/A _5620_/B _5634_/B vssd1 vssd1 vccd1 vccd1 _5979_/B sky130_fd_sc_hd__or3b_1
X_5551_ _5773_/A _6166_/A _5550_/Y vssd1 vssd1 vccd1 vccd1 _5556_/A sky130_fd_sc_hd__or3b_1
XFILLER_31_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8270_ _8450_/B _8270_/B vssd1 vssd1 vccd1 vccd1 _8463_/A sky130_fd_sc_hd__nand2_1
X_4502_ _5181_/A _4565_/B _5249_/A vssd1 vssd1 vccd1 vccd1 _4506_/B sky130_fd_sc_hd__o21ai_1
X_5482_ _5450_/X _5481_/Y _5478_/A _4616_/B vssd1 vssd1 vccd1 vccd1 _8712_/D sky130_fd_sc_hd__o2bb2a_1
X_7221_ _7221_/A _7221_/B vssd1 vssd1 vccd1 vccd1 _7221_/Y sky130_fd_sc_hd__nand2_1
X_4433_ _4457_/A vssd1 vssd1 vccd1 vccd1 _4438_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4364_ _4489_/A vssd1 vssd1 vccd1 vccd1 _4369_/A sky130_fd_sc_hd__clkbuf_2
X_7152_ _7515_/B _7518_/A _7515_/A vssd1 vssd1 vccd1 vccd1 _7516_/A sky130_fd_sc_hd__a21oi_1
X_6103_ _6103_/A _6163_/B vssd1 vssd1 vccd1 vccd1 _6104_/B sky130_fd_sc_hd__xnor2_2
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7083_ _7100_/A _7083_/B vssd1 vssd1 vccd1 vccd1 _7083_/Y sky130_fd_sc_hd__nand2_1
X_6034_ _6166_/A vssd1 vssd1 vccd1 vccd1 _6249_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_58_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7985_ _7919_/B _7919_/C _7919_/A vssd1 vssd1 vccd1 vccd1 _8004_/A sky130_fd_sc_hd__a21bo_1
XFILLER_54_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6936_ _6936_/A _6936_/B vssd1 vssd1 vccd1 vccd1 _6937_/B sky130_fd_sc_hd__xor2_1
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6867_ _7020_/B _6873_/A _6873_/B vssd1 vssd1 vccd1 vccd1 _6869_/B sky130_fd_sc_hd__or3_1
X_8606_ _8615_/A _8606_/B vssd1 vssd1 vccd1 vccd1 _8608_/A sky130_fd_sc_hd__or2_1
X_5818_ _5727_/A _5979_/B _5979_/C _6081_/A _5632_/A vssd1 vssd1 vccd1 vccd1 _5820_/B
+ sky130_fd_sc_hd__a32o_1
X_6798_ _6798_/A _7279_/A vssd1 vssd1 vccd1 vccd1 _7303_/A sky130_fd_sc_hd__nor2_4
X_8537_ _8537_/A _8537_/B vssd1 vssd1 vccd1 vccd1 _8538_/B sky130_fd_sc_hd__xnor2_1
X_5749_ _5749_/A _5837_/A vssd1 vssd1 vccd1 vccd1 _5754_/A sky130_fd_sc_hd__nor2_1
X_8468_ _8469_/A _8469_/B vssd1 vssd1 vccd1 vccd1 _8470_/A sky130_fd_sc_hd__and2_1
X_8399_ _8399_/A _8399_/B vssd1 vssd1 vccd1 vccd1 _8435_/B sky130_fd_sc_hd__xnor2_2
X_7419_ _7419_/A _7419_/B vssd1 vssd1 vccd1 vccd1 _7487_/A sky130_fd_sc_hd__xnor2_1
XFILLER_104_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7770_ _8182_/A _7836_/C _7882_/A _7882_/B vssd1 vssd1 vccd1 vccd1 _7772_/B sky130_fd_sc_hd__o22a_1
XFILLER_23_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4982_ _4982_/A _4982_/B vssd1 vssd1 vccd1 vccd1 _5005_/B sky130_fd_sc_hd__nor2_1
XFILLER_36_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6721_ _6721_/A _7137_/A vssd1 vssd1 vccd1 vccd1 _6722_/B sky130_fd_sc_hd__nand2_1
X_6652_ _7544_/A vssd1 vssd1 vccd1 vccd1 _7535_/A sky130_fd_sc_hd__clkinv_2
X_5603_ _5620_/A _5615_/B vssd1 vssd1 vccd1 vccd1 _5732_/A sky130_fd_sc_hd__or2_1
X_8322_ _8244_/A _8244_/B _8245_/B _8245_/A vssd1 vssd1 vccd1 vccd1 _8344_/A sky130_fd_sc_hd__o2bb2a_1
X_6583_ _6583_/A _6583_/B vssd1 vssd1 vccd1 vccd1 _6584_/B sky130_fd_sc_hd__nand2_1
X_5534_ _6378_/A _5533_/A _5861_/B _5533_/Y vssd1 vssd1 vccd1 vccd1 _5535_/B sky130_fd_sc_hd__o31a_1
XFILLER_11_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8253_ _8254_/A _8254_/B _8254_/C vssd1 vssd1 vccd1 vccd1 _8362_/A sky130_fd_sc_hd__o21ai_2
X_5465_ _5465_/A _5465_/B vssd1 vssd1 vccd1 vccd1 _5467_/A sky130_fd_sc_hd__nor2_1
X_4416_ _4419_/A vssd1 vssd1 vccd1 vccd1 _4416_/Y sky130_fd_sc_hd__inv_2
X_8184_ _8185_/A _8185_/B _8453_/A vssd1 vssd1 vccd1 vccd1 _8244_/A sky130_fd_sc_hd__a21oi_4
X_7204_ _7204_/A vssd1 vssd1 vccd1 vccd1 _7382_/A sky130_fd_sc_hd__clkbuf_2
X_7135_ _6809_/A _7078_/A _7105_/Y vssd1 vssd1 vccd1 vccd1 _7138_/B sky130_fd_sc_hd__a21oi_1
X_5396_ _8698_/Q _5394_/A _5392_/X vssd1 vssd1 vccd1 vccd1 _5397_/B sky130_fd_sc_hd__o21ai_1
XFILLER_101_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8860__77 vssd1 vssd1 vccd1 vccd1 _8860__77/HI _8969_/A sky130_fd_sc_hd__conb_1
X_7066_ _7067_/B _7067_/C _7067_/A vssd1 vssd1 vccd1 vccd1 _7068_/A sky130_fd_sc_hd__a21oi_1
X_6017_ _5861_/B _5913_/A _6016_/B vssd1 vssd1 vccd1 vccd1 _6017_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_39_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7968_ _7859_/A _7858_/B _7858_/A vssd1 vssd1 vccd1 vccd1 _7970_/B sky130_fd_sc_hd__o21ba_1
XFILLER_14_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7899_ _7899_/A vssd1 vssd1 vccd1 vccd1 _7996_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_52_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6919_ _7000_/B _6919_/B vssd1 vssd1 vccd1 vccd1 _6920_/B sky130_fd_sc_hd__and2_1
XFILLER_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5250_ _5263_/A _5250_/B _5250_/C _5250_/D vssd1 vssd1 vccd1 vccd1 _5250_/X sky130_fd_sc_hd__or4_1
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5181_ _5181_/A _5181_/B vssd1 vssd1 vccd1 vccd1 _5181_/Y sky130_fd_sc_hd__nand2_1
XFILLER_95_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8940_ _8940_/A _4429_/Y vssd1 vssd1 vccd1 vccd1 io_out[27] sky130_fd_sc_hd__ebufn_8
XFILLER_83_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7822_ _7915_/A vssd1 vssd1 vccd1 vccd1 _8568_/C sky130_fd_sc_hd__buf_2
XFILLER_64_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7753_ _7988_/A vssd1 vssd1 vccd1 vccd1 _8182_/A sky130_fd_sc_hd__clkbuf_2
X_4965_ _5209_/B _4995_/C _4964_/X vssd1 vssd1 vccd1 vccd1 _4965_/X sky130_fd_sc_hd__o21a_1
XFILLER_51_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6704_ _6704_/A _6704_/B vssd1 vssd1 vccd1 vccd1 _7034_/B sky130_fd_sc_hd__xnor2_4
X_7684_ _8771_/Q _7684_/B vssd1 vssd1 vccd1 vccd1 _7684_/X sky130_fd_sc_hd__and2b_1
X_4896_ _4912_/B _4922_/A vssd1 vssd1 vccd1 vccd1 _5087_/B sky130_fd_sc_hd__nor2_2
XFILLER_32_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6635_ _6635_/A vssd1 vssd1 vccd1 vccd1 _7141_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6566_ _6566_/A vssd1 vssd1 vccd1 vccd1 _8748_/D sky130_fd_sc_hd__clkbuf_1
X_8305_ _8305_/A _8305_/B vssd1 vssd1 vccd1 vccd1 _8306_/B sky130_fd_sc_hd__xnor2_1
X_5517_ _5505_/A _5505_/B _5508_/X _5509_/A vssd1 vssd1 vccd1 vccd1 _5521_/A sky130_fd_sc_hd__a31o_1
X_8236_ _8236_/A _8289_/B _8236_/C vssd1 vssd1 vccd1 vccd1 _8441_/A sky130_fd_sc_hd__or3_2
X_6497_ _8736_/Q _6497_/B _6497_/C vssd1 vssd1 vccd1 vccd1 _6501_/B sky130_fd_sc_hd__and3_1
X_5448_ _5448_/A vssd1 vssd1 vccd1 vccd1 _8707_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8167_ _8177_/A _8369_/A vssd1 vssd1 vccd1 vccd1 _8272_/D sky130_fd_sc_hd__nor2_1
X_5379_ _5381_/B _5379_/B _5389_/B vssd1 vssd1 vccd1 vccd1 _5380_/A sky130_fd_sc_hd__and3b_1
X_8098_ _8098_/A _8358_/A vssd1 vssd1 vccd1 vccd1 _8099_/D sky130_fd_sc_hd__or2b_1
X_7118_ _7118_/A _7118_/B vssd1 vssd1 vccd1 vccd1 _7123_/C sky130_fd_sc_hd__nor2_1
XFILLER_74_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7049_ _7120_/B _7049_/B vssd1 vssd1 vccd1 vccd1 _7221_/A sky130_fd_sc_hd__nor2_1
XFILLER_74_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4750_ _5300_/B _4751_/B vssd1 vssd1 vccd1 vccd1 _4752_/B sky130_fd_sc_hd__or2_1
X_4681_ _4807_/A vssd1 vssd1 vccd1 vccd1 _8588_/A sky130_fd_sc_hd__clkbuf_4
X_6420_ _6427_/B _6420_/B vssd1 vssd1 vccd1 vccd1 _6423_/C sky130_fd_sc_hd__and2b_1
X_6351_ _6351_/A _6351_/B vssd1 vssd1 vccd1 vccd1 _6351_/Y sky130_fd_sc_hd__nand2_1
X_5302_ _5302_/A _5302_/B vssd1 vssd1 vccd1 vccd1 _5302_/Y sky130_fd_sc_hd__nand2_1
X_6282_ _6326_/A _6326_/B vssd1 vssd1 vccd1 vccd1 _6283_/B sky130_fd_sc_hd__xor2_2
XFILLER_102_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8021_ _8059_/B _8020_/C _8020_/A vssd1 vssd1 vccd1 vccd1 _8039_/B sky130_fd_sc_hd__a21oi_2
X_5233_ _5215_/B _5142_/C _5211_/D _5197_/D vssd1 vssd1 vccd1 vccd1 _5234_/B sky130_fd_sc_hd__o31a_1
XFILLER_102_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5164_ _5164_/A _5201_/A vssd1 vssd1 vccd1 vccd1 _5164_/X sky130_fd_sc_hd__or2_1
XFILLER_56_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8830__47 vssd1 vssd1 vccd1 vccd1 _8830__47/HI _8939_/A sky130_fd_sc_hd__conb_1
XFILLER_96_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5095_ _5224_/B _5095_/B _5095_/C vssd1 vssd1 vccd1 vccd1 _5095_/X sky130_fd_sc_hd__or3_1
X_8923_ _8923_/A _4409_/Y vssd1 vssd1 vccd1 vccd1 io_out[10] sky130_fd_sc_hd__ebufn_8
XFILLER_17_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7805_ _8785_/Q _8661_/Q vssd1 vssd1 vccd1 vccd1 _8381_/A sky130_fd_sc_hd__and2b_2
X_5997_ _6088_/A _5998_/B vssd1 vssd1 vccd1 vccd1 _6075_/B sky130_fd_sc_hd__and2_1
X_8785_ _8785_/CLK _8785_/D vssd1 vssd1 vccd1 vccd1 _8785_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7736_ _7788_/A _7788_/B _7789_/B _7735_/X _7733_/A vssd1 vssd1 vccd1 vccd1 _7799_/B
+ sky130_fd_sc_hd__a311o_4
XFILLER_12_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4948_ _5159_/D _5054_/C vssd1 vssd1 vccd1 vccd1 _5209_/B sky130_fd_sc_hd__or2_2
X_7667_ _8628_/A _7667_/B vssd1 vssd1 vccd1 vccd1 _7667_/Y sky130_fd_sc_hd__nor2_1
X_4879_ _4902_/C _4879_/B vssd1 vssd1 vccd1 vccd1 _4879_/X sky130_fd_sc_hd__and2_1
XFILLER_20_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6618_ _6670_/A _6670_/B vssd1 vssd1 vccd1 vccd1 _7391_/A sky130_fd_sc_hd__xor2_4
X_7598_ _8615_/A vssd1 vssd1 vccd1 vccd1 _7598_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6549_ _8750_/Q vssd1 vssd1 vccd1 vccd1 _6628_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_8219_ _8220_/A _8220_/B vssd1 vssd1 vccd1 vccd1 _8221_/A sky130_fd_sc_hd__nand2_1
XFILLER_59_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5920_ _5920_/A _5920_/B vssd1 vssd1 vccd1 vccd1 _5922_/C sky130_fd_sc_hd__xnor2_1
XFILLER_80_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5851_ _5852_/A _6251_/A _5851_/C vssd1 vssd1 vccd1 vccd1 _5858_/B sky130_fd_sc_hd__and3_1
XFILLER_61_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5782_ _5783_/A _5783_/B vssd1 vssd1 vccd1 vccd1 _5872_/B sky130_fd_sc_hd__nor2_1
X_8570_ _8578_/A _8578_/B _8576_/B vssd1 vssd1 vccd1 vccd1 _8570_/X sky130_fd_sc_hd__or3_1
X_4802_ _4802_/A vssd1 vssd1 vccd1 vccd1 _8668_/D sky130_fd_sc_hd__clkbuf_1
X_7521_ _7521_/A _7523_/B vssd1 vssd1 vccd1 vccd1 _7522_/B sky130_fd_sc_hd__xnor2_1
X_4733_ _6613_/B _4733_/B _4733_/C vssd1 vssd1 vccd1 vccd1 _4973_/A sky130_fd_sc_hd__and3_1
X_7452_ _7390_/A _7390_/B _7451_/X vssd1 vssd1 vccd1 vccd1 _7453_/B sky130_fd_sc_hd__o21a_1
X_4664_ _4664_/A vssd1 vssd1 vccd1 vccd1 _8645_/D sky130_fd_sc_hd__clkbuf_1
X_6403_ _6403_/A vssd1 vssd1 vccd1 vccd1 _8718_/D sky130_fd_sc_hd__clkbuf_1
X_4595_ _8677_/Q _4595_/B vssd1 vssd1 vccd1 vccd1 _4596_/A sky130_fd_sc_hd__and2_2
X_7383_ _7383_/A _7383_/B vssd1 vssd1 vccd1 vccd1 _7384_/B sky130_fd_sc_hd__nor2_1
X_6334_ _6264_/A _6333_/Y _6180_/B vssd1 vssd1 vccd1 vccd1 _6334_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_103_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6265_ _6265_/A _6265_/B vssd1 vssd1 vccd1 vccd1 _6266_/B sky130_fd_sc_hd__xnor2_1
XFILLER_103_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8004_ _8004_/A _8061_/B _8004_/C vssd1 vssd1 vccd1 vccd1 _8060_/A sky130_fd_sc_hd__nand3_1
X_5216_ _5221_/A _5174_/A _5215_/X _5101_/B _4701_/A vssd1 vssd1 vccd1 vccd1 _5216_/X
+ sky130_fd_sc_hd__o32a_1
X_6196_ _6200_/A vssd1 vssd1 vccd1 vccd1 _6275_/S sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_84_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5147_ _5281_/B _5278_/B vssd1 vssd1 vccd1 vccd1 _5148_/C sky130_fd_sc_hd__nor2_1
XFILLER_28_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5078_ _5221_/C _5078_/B _5120_/B _5174_/B vssd1 vssd1 vccd1 vccd1 _5078_/X sky130_fd_sc_hd__or4_1
XFILLER_84_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8906_ _8906_/A _4388_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[25] sky130_fd_sc_hd__ebufn_8
X_8768_ _8771_/CLK _8768_/D vssd1 vssd1 vccd1 vccd1 _8768_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_12_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7719_ _7719_/A _7719_/B vssd1 vssd1 vccd1 vccd1 _7759_/A sky130_fd_sc_hd__xnor2_1
XFILLER_12_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8699_ _8732_/CLK _8699_/D vssd1 vssd1 vccd1 vccd1 _8699_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4380_ _4382_/A vssd1 vssd1 vccd1 vccd1 _4380_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6050_ _6050_/A _6050_/B vssd1 vssd1 vccd1 vccd1 _6050_/Y sky130_fd_sc_hd__nor2_1
XFILLER_98_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5001_ _5285_/A vssd1 vssd1 vccd1 vccd1 _5281_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_38_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8800__17 vssd1 vssd1 vccd1 vccd1 _8800__17/HI _8895_/A sky130_fd_sc_hd__conb_1
XFILLER_53_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6952_ _6994_/A _6994_/B vssd1 vssd1 vccd1 vccd1 _6953_/B sky130_fd_sc_hd__xnor2_1
XFILLER_38_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5903_ _5903_/A _5903_/B vssd1 vssd1 vccd1 vccd1 _5904_/B sky130_fd_sc_hd__or2_1
X_6883_ _6883_/A _6883_/B vssd1 vssd1 vccd1 vccd1 _6885_/A sky130_fd_sc_hd__xnor2_1
X_8622_ _8622_/A _8626_/B vssd1 vssd1 vccd1 vccd1 _8623_/B sky130_fd_sc_hd__nand2_1
X_5834_ _5980_/A vssd1 vssd1 vccd1 vccd1 _5897_/A sky130_fd_sc_hd__buf_2
XFILLER_22_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5765_ _5916_/B vssd1 vssd1 vccd1 vccd1 _5921_/B sky130_fd_sc_hd__clkbuf_2
X_8553_ _8562_/B _8562_/C _8562_/A vssd1 vssd1 vccd1 vccd1 _8563_/A sky130_fd_sc_hd__a21oi_1
X_5696_ _5805_/A _5805_/B vssd1 vssd1 vccd1 vccd1 _6398_/A sky130_fd_sc_hd__xnor2_1
X_8484_ _8550_/A _8484_/B vssd1 vssd1 vccd1 vccd1 _8549_/A sky130_fd_sc_hd__nand2_1
X_7504_ _7504_/A _7504_/B vssd1 vssd1 vccd1 vccd1 _7511_/A sky130_fd_sc_hd__xnor2_1
X_4716_ _4716_/A vssd1 vssd1 vccd1 vccd1 _5259_/D sky130_fd_sc_hd__clkbuf_2
X_4647_ _8640_/Q _4647_/B vssd1 vssd1 vccd1 vccd1 _4652_/C sky130_fd_sc_hd__and2_1
X_7435_ _7346_/A _7346_/B _7345_/B _7345_/A vssd1 vssd1 vccd1 vccd1 _7438_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7366_ _7366_/A _7508_/B vssd1 vssd1 vccd1 vccd1 _7367_/B sky130_fd_sc_hd__xnor2_1
X_6317_ _6257_/A _6257_/B _6256_/A vssd1 vssd1 vccd1 vccd1 _6318_/B sky130_fd_sc_hd__a21o_1
X_4578_ _8673_/Q _4584_/B vssd1 vssd1 vccd1 vccd1 _4579_/A sky130_fd_sc_hd__and2_1
X_7297_ _7209_/A _7297_/B vssd1 vssd1 vccd1 vccd1 _7297_/X sky130_fd_sc_hd__and2b_1
X_6248_ _6248_/A _6189_/B vssd1 vssd1 vccd1 vccd1 _6255_/B sky130_fd_sc_hd__or2b_1
X_6179_ _6101_/A _6207_/B _6100_/B _6102_/B _6102_/A vssd1 vssd1 vccd1 vccd1 _6244_/A
+ sky130_fd_sc_hd__a32oi_4
XFILLER_69_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8866__83 vssd1 vssd1 vccd1 vccd1 _8866__83/HI _8975_/A sky130_fd_sc_hd__conb_1
XFILLER_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5550_ _5916_/A _5527_/A _5662_/B _5549_/X vssd1 vssd1 vccd1 vccd1 _5550_/Y sky130_fd_sc_hd__a31oi_1
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4501_ _6655_/B vssd1 vssd1 vccd1 vccd1 _5249_/A sky130_fd_sc_hd__clkbuf_2
X_5481_ _5481_/A _5481_/B vssd1 vssd1 vccd1 vccd1 _5481_/Y sky130_fd_sc_hd__nand2_1
X_4432_ input1/X vssd1 vssd1 vccd1 vccd1 _4457_/A sky130_fd_sc_hd__clkbuf_2
X_7220_ _7220_/A _7220_/B vssd1 vssd1 vccd1 vccd1 _7240_/A sky130_fd_sc_hd__nor2_1
XFILLER_104_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7151_ _7151_/A _7151_/B vssd1 vssd1 vccd1 vccd1 _7515_/A sky130_fd_sc_hd__xnor2_1
X_4363_ _4363_/A vssd1 vssd1 vccd1 vccd1 _4363_/Y sky130_fd_sc_hd__inv_2
X_6102_ _6102_/A _6102_/B vssd1 vssd1 vccd1 vccd1 _6163_/B sky130_fd_sc_hd__xor2_2
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7082_ _7082_/A _7082_/B vssd1 vssd1 vccd1 vccd1 _7098_/B sky130_fd_sc_hd__xnor2_1
XFILLER_100_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6033_ _6238_/A _6106_/B vssd1 vssd1 vccd1 vccd1 _6036_/B sky130_fd_sc_hd__xor2_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7984_ _7930_/B _7930_/C _7930_/A vssd1 vssd1 vccd1 vccd1 _8016_/A sky130_fd_sc_hd__a21bo_1
XFILLER_26_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6935_ _6883_/A _6883_/B _6934_/X vssd1 vssd1 vccd1 vccd1 _6936_/B sky130_fd_sc_hd__o21a_1
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6866_ _6793_/C _6910_/A _6866_/C _6866_/D vssd1 vssd1 vccd1 vccd1 _6873_/B sky130_fd_sc_hd__and4b_1
XFILLER_34_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8605_ _8605_/A _8621_/B vssd1 vssd1 vccd1 vccd1 _8606_/B sky130_fd_sc_hd__nor2_1
X_5817_ _5837_/B vssd1 vssd1 vccd1 vccd1 _5986_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_22_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6797_ _6760_/X _6758_/Y _6759_/X _6752_/A vssd1 vssd1 vccd1 vccd1 _7279_/A sky130_fd_sc_hd__a31o_2
X_8536_ _8536_/A _8536_/B vssd1 vssd1 vccd1 vccd1 _8537_/B sky130_fd_sc_hd__xnor2_1
X_5748_ _5991_/A _5819_/C _5819_/D vssd1 vssd1 vccd1 vccd1 _5837_/A sky130_fd_sc_hd__or3_1
X_8467_ _8467_/A _8467_/B vssd1 vssd1 vccd1 vccd1 _8469_/B sky130_fd_sc_hd__xnor2_1
X_5679_ _5679_/A _5679_/B vssd1 vssd1 vccd1 vccd1 _5693_/A sky130_fd_sc_hd__nand2_1
X_8398_ _8396_/X _8398_/B vssd1 vssd1 vccd1 vccd1 _8399_/B sky130_fd_sc_hd__and2b_1
X_7418_ _7494_/A _7494_/B vssd1 vssd1 vccd1 vccd1 _7419_/B sky130_fd_sc_hd__xor2_1
XFILLER_89_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7349_ _7521_/A _7349_/B vssd1 vssd1 vccd1 vccd1 _7523_/A sky130_fd_sc_hd__and2_1
XFILLER_49_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4981_ _5040_/A _4883_/B _4982_/B vssd1 vssd1 vccd1 vccd1 _5269_/A sky130_fd_sc_hd__a21oi_2
X_6720_ _6721_/A _7137_/A vssd1 vssd1 vccd1 vccd1 _6729_/A sky130_fd_sc_hd__or2_1
X_6651_ _6651_/A _6651_/B vssd1 vssd1 vccd1 vccd1 _7544_/A sky130_fd_sc_hd__xnor2_2
X_5602_ _8723_/Q _8660_/Q vssd1 vssd1 vccd1 vccd1 _5615_/B sky130_fd_sc_hd__and2b_1
XFILLER_31_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6582_ _6583_/A _6588_/B vssd1 vssd1 vccd1 vccd1 _6582_/Y sky130_fd_sc_hd__nor2_1
X_8321_ _8306_/A _8306_/B _8320_/Y vssd1 vssd1 vccd1 vccd1 _8407_/B sky130_fd_sc_hd__a21o_1
X_5533_ _5533_/A _5683_/A vssd1 vssd1 vccd1 vccd1 _5533_/Y sky130_fd_sc_hd__nand2_1
XFILLER_8_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8252_ _8531_/A _8509_/A _8373_/A vssd1 vssd1 vccd1 vccd1 _8254_/C sky130_fd_sc_hd__o21a_1
X_5464_ _8710_/Q _5478_/B vssd1 vssd1 vccd1 vccd1 _5465_/B sky130_fd_sc_hd__and2b_1
X_4415_ _4419_/A vssd1 vssd1 vccd1 vccd1 _4415_/Y sky130_fd_sc_hd__inv_2
X_8183_ _8182_/B _8163_/B _8531_/A vssd1 vssd1 vccd1 vccd1 _8453_/A sky130_fd_sc_hd__a21o_2
X_7203_ _7301_/A _7370_/B vssd1 vssd1 vccd1 vccd1 _7208_/A sky130_fd_sc_hd__nand2_1
X_5395_ _8698_/Q _8697_/Q _5395_/C vssd1 vssd1 vccd1 vccd1 _5401_/C sky130_fd_sc_hd__and3_1
X_7134_ _7134_/A _7134_/B vssd1 vssd1 vccd1 vccd1 _7138_/A sky130_fd_sc_hd__xnor2_1
XFILLER_101_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7065_ _7346_/A _7065_/B vssd1 vssd1 vccd1 vccd1 _7067_/A sky130_fd_sc_hd__xnor2_1
X_6016_ _6016_/A _6016_/B vssd1 vssd1 vccd1 vccd1 _6019_/A sky130_fd_sc_hd__xnor2_1
XFILLER_100_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7967_ _7964_/X _7965_/Y _7892_/X _7893_/Y vssd1 vssd1 vccd1 vccd1 _7972_/B sky130_fd_sc_hd__o211a_1
XFILLER_42_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7898_ _7819_/A _7819_/B _7897_/X vssd1 vssd1 vccd1 vccd1 _7921_/A sky130_fd_sc_hd__a21o_1
X_6918_ _6918_/A _6918_/B vssd1 vssd1 vccd1 vccd1 _6919_/B sky130_fd_sc_hd__or2_1
XFILLER_42_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6849_ _7303_/A vssd1 vssd1 vccd1 vccd1 _7301_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_52_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8519_ _8519_/A _8519_/B vssd1 vssd1 vccd1 vccd1 _8535_/A sky130_fd_sc_hd__xnor2_1
XFILLER_2_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8836__53 vssd1 vssd1 vccd1 vccd1 _8836__53/HI _8945_/A sky130_fd_sc_hd__conb_1
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5180_ _5175_/X _5176_/X _5179_/X _5238_/B vssd1 vssd1 vccd1 vccd1 _5181_/B sky130_fd_sc_hd__o22ai_1
XFILLER_95_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7821_ _7821_/A _7821_/B vssd1 vssd1 vccd1 vccd1 _7915_/A sky130_fd_sc_hd__and2_1
XFILLER_64_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7752_ _7821_/A _7752_/B vssd1 vssd1 vccd1 vccd1 _7988_/A sky130_fd_sc_hd__xnor2_2
XFILLER_51_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4964_ _5145_/B vssd1 vssd1 vccd1 vccd1 _4964_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_51_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6703_ _6703_/A _6703_/B vssd1 vssd1 vccd1 vccd1 _6704_/B sky130_fd_sc_hd__nor2_2
X_7683_ _7671_/A _7708_/B _7678_/X _7676_/X vssd1 vssd1 vccd1 vccd1 _7688_/B sky130_fd_sc_hd__a211o_1
X_4895_ _5283_/B _5157_/A vssd1 vssd1 vccd1 vccd1 _5085_/A sky130_fd_sc_hd__or2_1
XFILLER_32_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6634_ _6793_/A _7198_/A vssd1 vssd1 vccd1 vccd1 _6635_/A sky130_fd_sc_hd__or2_1
X_6565_ _5389_/B _6568_/A _6621_/A vssd1 vssd1 vccd1 vccd1 _6566_/A sky130_fd_sc_hd__mux2_1
X_8304_ _8304_/A _8304_/B vssd1 vssd1 vccd1 vccd1 _8305_/B sky130_fd_sc_hd__nand2_1
X_5516_ _5852_/A _6142_/B vssd1 vssd1 vccd1 vccd1 _5533_/A sky130_fd_sc_hd__nand2_1
X_6496_ _6497_/B _6497_/C _6495_/Y vssd1 vssd1 vccd1 vccd1 _8735_/D sky130_fd_sc_hd__a21oi_1
X_8235_ _8206_/A _8206_/B _8234_/Y vssd1 vssd1 vccd1 vccd1 _8320_/A sky130_fd_sc_hd__a21oi_2
X_5447_ _5449_/A _5450_/A _5494_/A vssd1 vssd1 vccd1 vccd1 _5448_/A sky130_fd_sc_hd__mux2_1
X_8166_ _8270_/B _8389_/A _7755_/X vssd1 vssd1 vccd1 vccd1 _8369_/A sky130_fd_sc_hd__o21a_1
X_5378_ _6532_/D _5377_/C _8693_/Q vssd1 vssd1 vccd1 vccd1 _5379_/B sky130_fd_sc_hd__a21o_1
X_8097_ _8348_/A vssd1 vssd1 vccd1 vccd1 _8358_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7117_ _7117_/A _7117_/B vssd1 vssd1 vccd1 vccd1 _7130_/A sky130_fd_sc_hd__xnor2_1
X_7048_ _6922_/A _6922_/B _6938_/B _6939_/B _6939_/A vssd1 vssd1 vccd1 vccd1 _7163_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_101_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4680_ _4680_/A vssd1 vssd1 vccd1 vccd1 _8650_/D sky130_fd_sc_hd__clkbuf_1
X_6350_ _6016_/A _6252_/B _6251_/B vssd1 vssd1 vccd1 vccd1 _6353_/A sky130_fd_sc_hd__a21bo_1
X_5301_ _5301_/A _5301_/B _5301_/C _5300_/A vssd1 vssd1 vccd1 vccd1 _5302_/B sky130_fd_sc_hd__or4b_1
X_6281_ _6281_/A _6281_/B vssd1 vssd1 vccd1 vccd1 _6326_/B sky130_fd_sc_hd__xnor2_1
XFILLER_88_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8020_ _8020_/A _8059_/B _8020_/C vssd1 vssd1 vccd1 vccd1 _8058_/A sky130_fd_sc_hd__and3_1
X_5232_ _4697_/B _4702_/D _5225_/X _5231_/Y vssd1 vssd1 vccd1 vccd1 _5232_/X sky130_fd_sc_hd__o31a_1
X_5163_ _5163_/A _5163_/B _5163_/C vssd1 vssd1 vccd1 vccd1 _5265_/B sky130_fd_sc_hd__or3_2
XFILLER_68_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5094_ _5188_/B _5221_/C _5157_/B _4715_/B vssd1 vssd1 vccd1 vccd1 _5095_/B sky130_fd_sc_hd__o31a_1
X_8922_ _8922_/A _4407_/Y vssd1 vssd1 vccd1 vccd1 io_out[9] sky130_fd_sc_hd__ebufn_8
XFILLER_83_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7804_ _7804_/A vssd1 vssd1 vccd1 vccd1 _7813_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_24_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5996_ _5996_/A _6068_/C vssd1 vssd1 vccd1 vccd1 _5998_/B sky130_fd_sc_hd__xnor2_1
X_8784_ _8784_/CLK _8784_/D vssd1 vssd1 vccd1 vccd1 _8784_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_12_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7735_ _8605_/A _8658_/Q _8657_/Q _8599_/A vssd1 vssd1 vccd1 vccd1 _7735_/X sky130_fd_sc_hd__o211a_1
X_4947_ _4947_/A _4982_/B vssd1 vssd1 vccd1 vccd1 _5054_/C sky130_fd_sc_hd__nor2_1
XFILLER_24_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7666_ _7665_/X _7661_/A _7666_/S vssd1 vssd1 vccd1 vccd1 _7667_/B sky130_fd_sc_hd__mux2_1
XFILLER_32_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4878_ _4878_/A _4878_/B _4878_/C _4774_/A vssd1 vssd1 vccd1 vccd1 _4921_/A sky130_fd_sc_hd__or4b_2
X_6617_ _6617_/A _6617_/B vssd1 vssd1 vccd1 vccd1 _6670_/B sky130_fd_sc_hd__nor2_4
X_7597_ _8605_/A _8621_/B vssd1 vssd1 vccd1 vccd1 _8615_/A sky130_fd_sc_hd__and2_1
X_6548_ _8752_/Q vssd1 vssd1 vccd1 vccd1 _6593_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6479_ _8728_/Q _6452_/A _6473_/B _8730_/Q vssd1 vssd1 vccd1 vccd1 _6480_/B sky130_fd_sc_hd__a31o_1
X_8218_ _8304_/B _8218_/B vssd1 vssd1 vccd1 vccd1 _8220_/B sky130_fd_sc_hd__xnor2_1
XFILLER_87_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8149_ _8081_/B _8149_/B vssd1 vssd1 vccd1 vccd1 _8149_/X sky130_fd_sc_hd__and2b_1
X_8806__23 vssd1 vssd1 vccd1 vccd1 _8806__23/HI _8901_/A sky130_fd_sc_hd__conb_1
XINSDIODE2_0 _5076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5850_ _5913_/A vssd1 vssd1 vccd1 vccd1 _6251_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_61_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5781_ _5766_/C _5664_/B _5512_/B _5861_/B vssd1 vssd1 vccd1 vccd1 _5783_/B sky130_fd_sc_hd__o2bb2a_1
X_4801_ _7642_/A _4801_/B _4801_/C vssd1 vssd1 vccd1 vccd1 _4802_/A sky130_fd_sc_hd__and3_1
X_4732_ _4946_/A _4732_/B vssd1 vssd1 vccd1 vccd1 _4742_/A sky130_fd_sc_hd__nor2_1
XFILLER_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7520_ _7551_/A _7548_/A _7539_/A vssd1 vssd1 vccd1 vccd1 _7534_/A sky130_fd_sc_hd__a21oi_1
X_4663_ _4665_/B _4672_/B _4663_/C vssd1 vssd1 vccd1 vccd1 _4664_/A sky130_fd_sc_hd__and3b_1
X_7451_ _7451_/A _7394_/B vssd1 vssd1 vccd1 vccd1 _7451_/X sky130_fd_sc_hd__or2b_1
X_6402_ _5449_/A _5445_/A _6402_/S vssd1 vssd1 vccd1 vccd1 _6403_/A sky130_fd_sc_hd__mux2_1
X_4594_ _4594_/A vssd1 vssd1 vccd1 vccd1 _8930_/A sky130_fd_sc_hd__clkbuf_1
X_7382_ _7382_/A _7417_/B vssd1 vssd1 vccd1 vccd1 _7383_/B sky130_fd_sc_hd__and2_1
X_6333_ _6183_/A _5741_/A _5609_/Y vssd1 vssd1 vccd1 vccd1 _6333_/Y sky130_fd_sc_hd__o21ai_1
X_6264_ _6264_/A _6264_/B vssd1 vssd1 vccd1 vccd1 _6265_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8003_ _8061_/A _8002_/B _8002_/C vssd1 vssd1 vccd1 vccd1 _8004_/C sky130_fd_sc_hd__a21o_1
X_5215_ _5215_/A _5215_/B _5215_/C vssd1 vssd1 vccd1 vccd1 _5215_/X sky130_fd_sc_hd__or3_1
XFILLER_69_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6195_ _6259_/A _6259_/B vssd1 vssd1 vccd1 vccd1 _6260_/B sky130_fd_sc_hd__xor2_1
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5146_ _5201_/A vssd1 vssd1 vccd1 vccd1 _5278_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_84_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5077_ _5221_/B _5077_/B _5077_/C vssd1 vssd1 vccd1 vccd1 _5120_/B sky130_fd_sc_hd__or3_1
XFILLER_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8905_ _8905_/A _4387_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[24] sky130_fd_sc_hd__ebufn_8
XFILLER_25_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5979_ _5979_/A _5979_/B _5979_/C vssd1 vssd1 vccd1 vccd1 _5994_/B sky130_fd_sc_hd__and3_2
X_8767_ _8784_/CLK _8767_/D vssd1 vssd1 vccd1 vccd1 _8767_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7718_ _8568_/B _7706_/Y _8024_/A vssd1 vssd1 vccd1 vccd1 _7719_/B sky130_fd_sc_hd__o21a_1
XFILLER_100_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8698_ _8732_/CLK _8698_/D vssd1 vssd1 vccd1 vccd1 _8698_/Q sky130_fd_sc_hd__dfxtp_1
X_7649_ _7649_/A _7649_/B vssd1 vssd1 vccd1 vccd1 _7649_/X sky130_fd_sc_hd__or2_1
XFILLER_79_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5000_ _5123_/A vssd1 vssd1 vccd1 vccd1 _5285_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8797__14 vssd1 vssd1 vccd1 vccd1 _8797__14/HI _8892_/A sky130_fd_sc_hd__conb_1
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6951_ _7373_/A _7047_/B vssd1 vssd1 vccd1 vccd1 _6994_/B sky130_fd_sc_hd__xnor2_1
X_5902_ _5903_/A _5903_/B vssd1 vssd1 vccd1 vccd1 _6007_/B sky130_fd_sc_hd__nand2_1
X_6882_ _7380_/A _7311_/S vssd1 vssd1 vccd1 vccd1 _6883_/B sky130_fd_sc_hd__xnor2_1
XFILLER_46_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5833_ _5889_/B _5832_/C _5832_/A vssd1 vssd1 vccd1 vccd1 _5841_/B sky130_fd_sc_hd__a21o_1
X_8621_ _8784_/Q _8621_/B vssd1 vssd1 vccd1 vccd1 _8626_/B sky130_fd_sc_hd__or2_1
X_8552_ _8552_/A _8552_/B vssd1 vssd1 vccd1 vccd1 _8554_/A sky130_fd_sc_hd__xor2_1
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5764_ _5764_/A _5764_/B vssd1 vssd1 vccd1 vccd1 _5864_/A sky130_fd_sc_hd__nor2_1
X_7503_ _7503_/A _7503_/B vssd1 vssd1 vccd1 vccd1 _7504_/B sky130_fd_sc_hd__xnor2_1
X_5695_ _5681_/A _6378_/B _5697_/B _5694_/A vssd1 vssd1 vccd1 vccd1 _5805_/B sky130_fd_sc_hd__a31o_1
X_8483_ _8483_/A _8483_/B vssd1 vssd1 vccd1 vccd1 _8484_/B sky130_fd_sc_hd__or2_1
X_4715_ _5182_/A _4715_/B vssd1 vssd1 vccd1 vccd1 _4716_/A sky130_fd_sc_hd__nor2_4
X_7434_ _7434_/A _7434_/B vssd1 vssd1 vccd1 vccd1 _7438_/A sky130_fd_sc_hd__xnor2_2
X_4646_ _4646_/A vssd1 vssd1 vccd1 vccd1 _8639_/D sky130_fd_sc_hd__clkbuf_1
X_4577_ _4577_/A vssd1 vssd1 vccd1 vccd1 _8926_/A sky130_fd_sc_hd__clkbuf_1
X_7365_ _7389_/A _6816_/A _7312_/B _7228_/A vssd1 vssd1 vccd1 vccd1 _7508_/B sky130_fd_sc_hd__a22oi_4
XFILLER_30_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6316_ _6316_/A _6316_/B vssd1 vssd1 vccd1 vccd1 _6355_/A sky130_fd_sc_hd__xnor2_1
X_7296_ _7427_/A _7427_/B vssd1 vssd1 vccd1 vccd1 _7321_/A sky130_fd_sc_hd__xnor2_2
XFILLER_39_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6247_ _6247_/A _6188_/A vssd1 vssd1 vccd1 vccd1 _6255_/A sky130_fd_sc_hd__or2b_1
X_6178_ _6178_/A _6178_/B vssd1 vssd1 vccd1 vccd1 _6243_/A sky130_fd_sc_hd__xnor2_1
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5129_ _5150_/A _5122_/Y _5128_/Y _4819_/A vssd1 vssd1 vccd1 vccd1 _5129_/X sky130_fd_sc_hd__a211o_1
XFILLER_84_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4500_ _8659_/Q vssd1 vssd1 vccd1 vccd1 _6655_/B sky130_fd_sc_hd__buf_2
X_5480_ _5480_/A _5485_/S _5480_/C _5484_/B vssd1 vssd1 vccd1 vccd1 _5481_/B sky130_fd_sc_hd__nand4_1
X_4431_ _4431_/A vssd1 vssd1 vccd1 vccd1 _4431_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7150_ _7538_/A _7537_/A vssd1 vssd1 vccd1 vccd1 _7518_/A sky130_fd_sc_hd__nand2_1
X_4362_ _4363_/A vssd1 vssd1 vccd1 vccd1 _4362_/Y sky130_fd_sc_hd__inv_2
X_6101_ _6101_/A _6101_/B vssd1 vssd1 vccd1 vccd1 _6102_/B sky130_fd_sc_hd__xnor2_2
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7081_ _7087_/A _7087_/B vssd1 vssd1 vccd1 vccd1 _7082_/B sky130_fd_sc_hd__xor2_1
X_6032_ _5920_/A _5918_/X _6171_/A _5856_/A vssd1 vssd1 vccd1 vccd1 _6106_/B sky130_fd_sc_hd__o22ai_2
XFILLER_86_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7983_ _7934_/A _7934_/B _7934_/D _7982_/X vssd1 vssd1 vccd1 vccd1 _8020_/A sky130_fd_sc_hd__a31o_1
X_6934_ _6886_/A _7303_/A _6883_/A _6883_/B vssd1 vssd1 vccd1 vccd1 _6934_/X sky130_fd_sc_hd__a22o_1
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8604_ _7734_/A _7627_/X _8603_/X _7642_/X vssd1 vssd1 vccd1 vccd1 _8781_/D sky130_fd_sc_hd__o211a_1
XFILLER_62_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6865_ _6765_/A _6836_/A _6910_/A _6910_/B _6866_/C vssd1 vssd1 vccd1 vccd1 _6873_/A
+ sky130_fd_sc_hd__a32oi_4
X_5816_ _5891_/A _5983_/A vssd1 vssd1 vccd1 vccd1 _5837_/B sky130_fd_sc_hd__nor2_1
X_6796_ _6960_/B _7123_/B vssd1 vssd1 vccd1 vccd1 _6801_/A sky130_fd_sc_hd__nand2_1
X_8535_ _8535_/A _8535_/B vssd1 vssd1 vccd1 vccd1 _8536_/B sky130_fd_sc_hd__xnor2_1
X_5747_ _5746_/B _5746_/C _5746_/A vssd1 vssd1 vccd1 vccd1 _5756_/B sky130_fd_sc_hd__a21o_1
X_8466_ _8521_/A _8521_/B vssd1 vssd1 vccd1 vccd1 _8467_/B sky130_fd_sc_hd__xnor2_1
X_5678_ _5678_/A _5678_/B vssd1 vssd1 vccd1 vccd1 _5679_/B sky130_fd_sc_hd__nand2_1
X_7417_ _7417_/A _7417_/B vssd1 vssd1 vccd1 vccd1 _7494_/B sky130_fd_sc_hd__xnor2_2
X_8397_ _8396_/B _8396_/C _8396_/A vssd1 vssd1 vccd1 vccd1 _8398_/B sky130_fd_sc_hd__a21o_1
X_4629_ _8634_/Q _4631_/C _4628_/X vssd1 vssd1 vccd1 vccd1 _4630_/B sky130_fd_sc_hd__o21ai_1
X_7348_ _7348_/A _7348_/B _7348_/C vssd1 vssd1 vccd1 vccd1 _7349_/B sky130_fd_sc_hd__nand3_1
XFILLER_1_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7279_ _7279_/A _7279_/B vssd1 vssd1 vccd1 vccd1 _7281_/A sky130_fd_sc_hd__nor2_1
XFILLER_89_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4980_ _5271_/A _5149_/C _4980_/C _5096_/B vssd1 vssd1 vccd1 vccd1 _4980_/X sky130_fd_sc_hd__or4_1
XFILLER_63_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6650_ _6650_/A _6924_/A vssd1 vssd1 vccd1 vccd1 _6651_/B sky130_fd_sc_hd__nor2_1
XFILLER_31_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5601_ _8660_/Q _8723_/Q vssd1 vssd1 vccd1 vccd1 _5620_/A sky130_fd_sc_hd__and2b_1
X_6581_ _6628_/B _6567_/X _6569_/X _6580_/X vssd1 vssd1 vccd1 vccd1 _8750_/D sky130_fd_sc_hd__a22o_1
X_8320_ _8320_/A _8320_/B vssd1 vssd1 vccd1 vccd1 _8320_/Y sky130_fd_sc_hd__nor2_1
X_5532_ _5532_/A _5531_/X vssd1 vssd1 vccd1 vccd1 _5683_/A sky130_fd_sc_hd__or2b_1
X_8251_ _8439_/A _8531_/A vssd1 vssd1 vccd1 vccd1 _8373_/A sky130_fd_sc_hd__nand2_1
X_5463_ _5477_/B _5463_/B vssd1 vssd1 vccd1 vccd1 _5465_/A sky130_fd_sc_hd__and2b_1
X_4414_ _4426_/A vssd1 vssd1 vccd1 vccd1 _4419_/A sky130_fd_sc_hd__buf_2
XFILLER_99_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8182_ _8182_/A _8182_/B vssd1 vssd1 vccd1 vccd1 _8531_/A sky130_fd_sc_hd__nor2_2
X_7202_ _7331_/A vssd1 vssd1 vccd1 vccd1 _7370_/B sky130_fd_sc_hd__clkbuf_2
X_5394_ _5394_/A _5394_/B vssd1 vssd1 vccd1 vccd1 _8697_/D sky130_fd_sc_hd__nor2_1
X_7133_ _7154_/B _7133_/B vssd1 vssd1 vccd1 vccd1 _7519_/A sky130_fd_sc_hd__xnor2_1
XFILLER_98_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7064_ _7064_/A _7064_/B vssd1 vssd1 vccd1 vccd1 _7065_/B sky130_fd_sc_hd__xor2_1
XFILLER_100_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6015_ _6059_/A _6228_/A _6014_/Y vssd1 vssd1 vccd1 vccd1 _6016_/B sky130_fd_sc_hd__o21bai_2
XFILLER_39_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7966_ _7892_/X _7893_/Y _7964_/X _7965_/Y vssd1 vssd1 vccd1 vccd1 _7972_/A sky130_fd_sc_hd__a211oi_2
XFILLER_54_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7897_ _8450_/B _7897_/B vssd1 vssd1 vccd1 vccd1 _7897_/X sky130_fd_sc_hd__and2_1
X_6917_ _6918_/A _6918_/B vssd1 vssd1 vccd1 vccd1 _7000_/B sky130_fd_sc_hd__nand2_1
X_6848_ _6848_/A _6848_/B vssd1 vssd1 vccd1 vccd1 _6894_/A sky130_fd_sc_hd__nand2_1
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8518_ _8518_/A _8518_/B vssd1 vssd1 vccd1 vccd1 _8519_/B sky130_fd_sc_hd__nor2_1
XFILLER_10_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6779_ _6960_/B _6779_/B vssd1 vssd1 vccd1 vccd1 _6840_/A sky130_fd_sc_hd__xor2_1
X_8449_ _8163_/A _8165_/B _8261_/A vssd1 vssd1 vccd1 vccd1 _8449_/X sky130_fd_sc_hd__a21o_1
XFILLER_2_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8851__68 vssd1 vssd1 vccd1 vccd1 _8851__68/HI _8960_/A sky130_fd_sc_hd__conb_1
XFILLER_58_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7820_ _7820_/A _7895_/C vssd1 vssd1 vccd1 vccd1 _7831_/A sky130_fd_sc_hd__xnor2_1
XFILLER_64_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7751_ _7934_/A _8450_/B vssd1 vssd1 vccd1 vccd1 _7836_/C sky130_fd_sc_hd__nand2_1
XFILLER_51_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4963_ _5042_/A vssd1 vssd1 vccd1 vccd1 _5145_/B sky130_fd_sc_hd__buf_2
X_7682_ _7693_/A vssd1 vssd1 vccd1 vccd1 _8024_/A sky130_fd_sc_hd__inv_2
X_6702_ _6702_/A vssd1 vssd1 vccd1 vccd1 _6703_/A sky130_fd_sc_hd__inv_2
X_4894_ _4910_/A _4894_/B vssd1 vssd1 vccd1 vccd1 _5157_/A sky130_fd_sc_hd__nor2_1
X_6633_ _6898_/A _6774_/A vssd1 vssd1 vccd1 vccd1 _7198_/A sky130_fd_sc_hd__or2_2
XFILLER_32_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6564_ _8748_/Q vssd1 vssd1 vccd1 vccd1 _6621_/A sky130_fd_sc_hd__inv_2
X_8303_ _8303_/A _8303_/B vssd1 vssd1 vccd1 vccd1 _8305_/A sky130_fd_sc_hd__nor2_1
X_5515_ _5853_/A vssd1 vssd1 vccd1 vccd1 _6142_/B sky130_fd_sc_hd__clkbuf_2
X_6495_ _6497_/B _6497_/C _6524_/B vssd1 vssd1 vccd1 vccd1 _6495_/Y sky130_fd_sc_hd__o21ai_1
X_8234_ _8234_/A _8234_/B vssd1 vssd1 vccd1 vccd1 _8234_/Y sky130_fd_sc_hd__nor2_1
X_5446_ _8707_/Q vssd1 vssd1 vccd1 vccd1 _5494_/A sky130_fd_sc_hd__inv_2
XFILLER_87_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8165_ _8273_/B _8165_/B _8165_/C vssd1 vssd1 vccd1 vccd1 _8389_/A sky130_fd_sc_hd__and3b_1
X_5377_ _8693_/Q _8692_/Q _5377_/C vssd1 vssd1 vccd1 vccd1 _5381_/B sky130_fd_sc_hd__and3_1
XFILLER_101_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8096_ _8198_/A _8096_/B vssd1 vssd1 vccd1 vccd1 _8099_/C sky130_fd_sc_hd__xnor2_1
XFILLER_59_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7116_ _7116_/A _7116_/B vssd1 vssd1 vccd1 vccd1 _7154_/B sky130_fd_sc_hd__xnor2_1
XFILLER_101_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7047_ _7484_/S _7047_/B vssd1 vssd1 vccd1 vccd1 _7060_/A sky130_fd_sc_hd__and2_1
XFILLER_86_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7949_ _8044_/A _7949_/B vssd1 vssd1 vccd1 vccd1 _8023_/B sky130_fd_sc_hd__nor2_2
XFILLER_15_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5300_ _5300_/A _5300_/B _5300_/C _5301_/A vssd1 vssd1 vccd1 vccd1 _5302_/A sky130_fd_sc_hd__or4b_1
X_6280_ _6280_/A _6280_/B vssd1 vssd1 vccd1 vccd1 _6281_/B sky130_fd_sc_hd__xor2_1
XFILLER_69_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5231_ _5231_/A _5231_/B vssd1 vssd1 vccd1 vccd1 _5231_/Y sky130_fd_sc_hd__nand2_1
X_5162_ _5162_/A vssd1 vssd1 vccd1 vccd1 _5278_/A sky130_fd_sc_hd__inv_2
X_5093_ _5227_/A _5078_/X _5084_/X _5092_/X vssd1 vssd1 vccd1 vccd1 _5093_/X sky130_fd_sc_hd__o31a_1
XFILLER_68_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8921_ _8921_/A _4406_/Y vssd1 vssd1 vccd1 vccd1 io_out[8] sky130_fd_sc_hd__ebufn_8
XFILLER_83_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7803_ _8163_/A _7897_/B vssd1 vssd1 vccd1 vccd1 _7819_/A sky130_fd_sc_hd__xnor2_1
X_8783_ _8783_/CLK _8783_/D vssd1 vssd1 vccd1 vccd1 _8783_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7734_ _7734_/A vssd1 vssd1 vccd1 vccd1 _8599_/A sky130_fd_sc_hd__inv_2
X_5995_ _5995_/A _5995_/B vssd1 vssd1 vccd1 vccd1 _6068_/C sky130_fd_sc_hd__xor2_1
XFILLER_52_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4946_ _4946_/A _5174_/A _4995_/C vssd1 vssd1 vccd1 vccd1 _4946_/X sky130_fd_sc_hd__or3_1
X_7665_ _7665_/A _7665_/B vssd1 vssd1 vccd1 vccd1 _7665_/X sky130_fd_sc_hd__or2_1
X_4877_ _4877_/A _4877_/B _4877_/C vssd1 vssd1 vccd1 vccd1 _4922_/A sky130_fd_sc_hd__or3_2
X_7596_ _8612_/B vssd1 vssd1 vccd1 vccd1 _8621_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6616_ _6615_/B _8761_/Q vssd1 vssd1 vccd1 vccd1 _6617_/B sky130_fd_sc_hd__and2b_1
X_6547_ _6537_/X _6546_/Y _7621_/A vssd1 vssd1 vccd1 vccd1 _8746_/D sky130_fd_sc_hd__o21a_1
X_6478_ _8729_/Q _8730_/Q _6478_/C vssd1 vssd1 vccd1 vccd1 _6486_/C sky130_fd_sc_hd__and3_1
X_8217_ _8124_/A _8124_/C _8124_/B vssd1 vssd1 vccd1 vccd1 _8218_/B sky130_fd_sc_hd__a21boi_1
X_5429_ _5429_/A vssd1 vssd1 vccd1 vccd1 _8705_/D sky130_fd_sc_hd__clkinv_2
X_8148_ _8117_/A _8117_/B _8147_/Y vssd1 vssd1 vccd1 vccd1 _8232_/A sky130_fd_sc_hd__a21boi_2
XFILLER_59_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_1 _5280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8821__38 vssd1 vssd1 vccd1 vccd1 _8821__38/HI _8916_/A sky130_fd_sc_hd__conb_1
X_8079_ _8185_/B _8079_/B vssd1 vssd1 vccd1 vccd1 _8080_/B sky130_fd_sc_hd__nand2_1
XFILLER_74_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_0_0_wb_clk_i clkbuf_4_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _8704_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_19_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4800_ _4804_/B _4804_/C vssd1 vssd1 vccd1 vccd1 _4801_/C sky130_fd_sc_hd__nand2_1
X_5780_ _5864_/A _5864_/B vssd1 vssd1 vccd1 vccd1 _5786_/A sky130_fd_sc_hd__xnor2_1
XFILLER_34_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4731_ _5271_/A _4730_/A _4730_/Y _4705_/X vssd1 vssd1 vccd1 vccd1 _8655_/D sky130_fd_sc_hd__o211a_1
XFILLER_21_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4662_ _8644_/Q _8643_/Q _4656_/B _8645_/Q vssd1 vssd1 vccd1 vccd1 _4663_/C sky130_fd_sc_hd__a31o_1
X_7450_ _7388_/S _7391_/Y _7450_/S vssd1 vssd1 vccd1 vccd1 _7453_/A sky130_fd_sc_hd__mux2_1
X_6401_ _6387_/X _6383_/X _6399_/X _6400_/Y vssd1 vssd1 vccd1 vccd1 _8717_/D sky130_fd_sc_hd__a31oi_1
X_4593_ _8676_/Q _4595_/B vssd1 vssd1 vccd1 vccd1 _4594_/A sky130_fd_sc_hd__and2_1
X_7381_ _7382_/A _7417_/B vssd1 vssd1 vccd1 vccd1 _7383_/A sky130_fd_sc_hd__nor2_1
X_6332_ _6271_/A _6271_/B _6269_/A vssd1 vssd1 vccd1 vccd1 _6336_/A sky130_fd_sc_hd__o21a_1
X_6263_ _6263_/A _6263_/B vssd1 vssd1 vccd1 vccd1 _6264_/B sky130_fd_sc_hd__xnor2_1
X_8002_ _8061_/A _8002_/B _8002_/C vssd1 vssd1 vccd1 vccd1 _8061_/B sky130_fd_sc_hd__nand3_1
X_5214_ _5047_/A _5221_/C _5207_/B _5031_/B vssd1 vssd1 vccd1 vccd1 _5214_/X sky130_fd_sc_hd__o31a_1
X_6194_ _6194_/A _6194_/B vssd1 vssd1 vccd1 vccd1 _6259_/B sky130_fd_sc_hd__xor2_1
XFILLER_96_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5145_ _5168_/A _5145_/B vssd1 vssd1 vccd1 vccd1 _5145_/Y sky130_fd_sc_hd__nor2_1
XFILLER_56_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5076_ _5076_/A vssd1 vssd1 vccd1 vccd1 _5221_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_8904_ _8904_/A _4386_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[23] sky130_fd_sc_hd__ebufn_8
XFILLER_25_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5978_ _6004_/B _5897_/B _5977_/Y vssd1 vssd1 vccd1 vccd1 _6077_/A sky130_fd_sc_hd__a21bo_1
XFILLER_52_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8766_ _8784_/CLK _8766_/D vssd1 vssd1 vccd1 vccd1 _8766_/Q sky130_fd_sc_hd__dfxtp_1
X_7717_ _7839_/B vssd1 vssd1 vccd1 vccd1 _8568_/B sky130_fd_sc_hd__clkbuf_2
X_4929_ _5076_/A _5171_/B vssd1 vssd1 vccd1 vccd1 _5136_/B sky130_fd_sc_hd__or2_2
X_8697_ _8704_/CLK _8697_/D vssd1 vssd1 vccd1 vccd1 _8697_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7648_ _7652_/B _7648_/B vssd1 vssd1 vccd1 vccd1 _7648_/Y sky130_fd_sc_hd__nor2_1
XFILLER_20_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7579_ _7583_/A _7579_/B vssd1 vssd1 vccd1 vccd1 _7579_/Y sky130_fd_sc_hd__nand2_1
XFILLER_4_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6950_ _6816_/A _6948_/Y _7049_/B _6818_/A vssd1 vssd1 vccd1 vccd1 _7047_/B sky130_fd_sc_hd__a31o_1
XFILLER_19_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5901_ _5977_/B _6002_/A vssd1 vssd1 vccd1 vccd1 _5903_/B sky130_fd_sc_hd__xnor2_1
XFILLER_19_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6881_ _6881_/A _6881_/B vssd1 vssd1 vccd1 vccd1 _6887_/A sky130_fd_sc_hd__nand2_1
X_5832_ _5832_/A _5889_/B _5832_/C vssd1 vssd1 vccd1 vccd1 _5888_/A sky130_fd_sc_hd__nand3_1
X_8620_ _8784_/Q _8621_/B vssd1 vssd1 vccd1 vccd1 _8622_/A sky130_fd_sc_hd__nand2_1
X_5763_ _5810_/B _5810_/C _5810_/A vssd1 vssd1 vccd1 vccd1 _5792_/B sky130_fd_sc_hd__a21o_1
X_8551_ _8548_/Y _8549_/X _8550_/X vssd1 vssd1 vccd1 vccd1 _8565_/C sky130_fd_sc_hd__o21ai_1
X_7502_ _7502_/A _7502_/B vssd1 vssd1 vccd1 vccd1 _7503_/B sky130_fd_sc_hd__xnor2_1
X_4714_ _5042_/A vssd1 vssd1 vccd1 vccd1 _4715_/B sky130_fd_sc_hd__buf_2
X_5694_ _5694_/A _5694_/B vssd1 vssd1 vccd1 vccd1 _5697_/B sky130_fd_sc_hd__nor2_1
X_8482_ _8483_/A _8483_/B vssd1 vssd1 vccd1 vccd1 _8550_/A sky130_fd_sc_hd__nand2_1
X_7433_ _7433_/A _7433_/B vssd1 vssd1 vccd1 vccd1 _7434_/B sky130_fd_sc_hd__xnor2_2
X_4645_ _4647_/B _4672_/B _4645_/C vssd1 vssd1 vccd1 vccd1 _4646_/A sky130_fd_sc_hd__and3b_1
X_4576_ _8672_/Q _4584_/B vssd1 vssd1 vccd1 vccd1 _4577_/A sky130_fd_sc_hd__and2_1
X_7364_ _7460_/S _7227_/A _7370_/B _7331_/B vssd1 vssd1 vccd1 vccd1 _7367_/A sky130_fd_sc_hd__a22o_1
X_6315_ _6315_/A _6315_/B vssd1 vssd1 vccd1 vccd1 _6316_/B sky130_fd_sc_hd__xnor2_1
XFILLER_89_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7295_ _7318_/B _7180_/B _7194_/B _7294_/Y vssd1 vssd1 vccd1 vccd1 _7427_/B sky130_fd_sc_hd__a31o_1
XFILLER_103_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6246_ _6252_/A _6246_/B vssd1 vssd1 vccd1 vccd1 _6257_/A sky130_fd_sc_hd__nor2_1
XFILLER_103_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6177_ _6177_/A _6177_/B vssd1 vssd1 vccd1 vccd1 _6178_/B sky130_fd_sc_hd__xor2_1
XFILLER_69_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5128_ _5128_/A _5128_/B vssd1 vssd1 vccd1 vccd1 _5128_/Y sky130_fd_sc_hd__nor2_1
XFILLER_72_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5059_ _5201_/A _5059_/B vssd1 vssd1 vccd1 vccd1 _5274_/B sky130_fd_sc_hd__or2_2
XFILLER_13_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8749_ _8753_/CLK _8749_/D vssd1 vssd1 vccd1 vccd1 _8749_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4430_ _4431_/A vssd1 vssd1 vccd1 vccd1 _4430_/Y sky130_fd_sc_hd__inv_2
X_8857__74 vssd1 vssd1 vccd1 vccd1 _8857__74/HI _8966_/A sky130_fd_sc_hd__conb_1
XFILLER_6_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6100_ _6207_/B _6100_/B vssd1 vssd1 vccd1 vccd1 _6101_/B sky130_fd_sc_hd__nand2_1
XFILLER_6_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4361_ _4363_/A vssd1 vssd1 vccd1 vccd1 _4361_/Y sky130_fd_sc_hd__inv_2
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7080_ _7141_/A _7400_/B _7080_/C _7080_/D vssd1 vssd1 vccd1 vccd1 _7087_/B sky130_fd_sc_hd__or4_2
X_6031_ _5938_/A _5938_/B _5939_/A vssd1 vssd1 vccd1 vccd1 _6042_/A sky130_fd_sc_hd__a21oi_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7982_ _7982_/A _7982_/B _7982_/C vssd1 vssd1 vccd1 vccd1 _7982_/X sky130_fd_sc_hd__and3_1
XFILLER_54_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6933_ _6933_/A _6933_/B vssd1 vssd1 vccd1 vccd1 _6936_/A sky130_fd_sc_hd__xnor2_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6864_ _6769_/A _6837_/B _6862_/X _6876_/A vssd1 vssd1 vccd1 vccd1 _6883_/A sky130_fd_sc_hd__a31o_2
XFILLER_34_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5815_ _5835_/A _5728_/B _5728_/C vssd1 vssd1 vccd1 vccd1 _5822_/A sky130_fd_sc_hd__o21bai_1
X_8603_ _8603_/A _8603_/B vssd1 vssd1 vccd1 vccd1 _8603_/X sky130_fd_sc_hd__or2_1
XFILLER_50_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6795_ _6863_/C vssd1 vssd1 vccd1 vccd1 _7123_/B sky130_fd_sc_hd__buf_2
X_8534_ _8534_/A _8534_/B vssd1 vssd1 vccd1 vccd1 _8535_/B sky130_fd_sc_hd__xnor2_1
X_5746_ _5746_/A _5746_/B _5746_/C vssd1 vssd1 vccd1 vccd1 _5756_/A sky130_fd_sc_hd__nand3_1
XFILLER_22_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8465_ _8465_/A _8465_/B vssd1 vssd1 vccd1 vccd1 _8521_/B sky130_fd_sc_hd__xnor2_1
X_5677_ _5677_/A _5677_/B vssd1 vssd1 vccd1 vccd1 _5805_/A sky130_fd_sc_hd__xor2_1
X_4628_ _4672_/B vssd1 vssd1 vccd1 vccd1 _4628_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7416_ _7416_/A _7416_/B vssd1 vssd1 vccd1 vccd1 _7494_/A sky130_fd_sc_hd__nor2_1
X_8396_ _8396_/A _8396_/B _8396_/C vssd1 vssd1 vccd1 vccd1 _8396_/X sky130_fd_sc_hd__and3_1
XFILLER_104_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7347_ _7348_/A _7348_/B _7348_/C vssd1 vssd1 vccd1 vccd1 _7521_/A sky130_fd_sc_hd__a21o_1
X_4559_ _8653_/Q vssd1 vssd1 vccd1 vccd1 _5138_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_103_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7278_ _7278_/A _7278_/B vssd1 vssd1 vccd1 vccd1 _7293_/A sky130_fd_sc_hd__nor2_1
XFILLER_103_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6229_ _6228_/Y _6168_/B _6166_/X vssd1 vssd1 vccd1 vccd1 _6231_/A sky130_fd_sc_hd__a21boi_1
XFILLER_66_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5600_ _6068_/A _6004_/A vssd1 vssd1 vccd1 vccd1 _5628_/A sky130_fd_sc_hd__nand2_1
X_6580_ _6580_/A _6580_/B vssd1 vssd1 vccd1 vccd1 _6580_/X sky130_fd_sc_hd__xor2_1
X_5531_ _5773_/A _5682_/B _6142_/B _5531_/D vssd1 vssd1 vccd1 vccd1 _5531_/X sky130_fd_sc_hd__or4_1
X_8250_ _8371_/A _8568_/C _8389_/B vssd1 vssd1 vccd1 vccd1 _8509_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5462_ _5462_/A _5462_/B vssd1 vssd1 vccd1 vccd1 _5462_/X sky130_fd_sc_hd__and2_1
X_7201_ _7038_/A _7038_/B _7200_/X vssd1 vssd1 vccd1 vccd1 _7209_/A sky130_fd_sc_hd__a21oi_1
X_4413_ _4413_/A vssd1 vssd1 vccd1 vccd1 _4413_/Y sky130_fd_sc_hd__clkinv_2
X_8181_ _8181_/A _8181_/B vssd1 vssd1 vccd1 vccd1 _8185_/A sky130_fd_sc_hd__or2_1
X_5393_ _8697_/Q _5395_/C _5392_/X vssd1 vssd1 vccd1 vccd1 _5394_/B sky130_fd_sc_hd__o21ai_1
X_7132_ _7137_/A _7137_/B _7131_/X vssd1 vssd1 vccd1 vccd1 _7133_/B sky130_fd_sc_hd__o21a_1
XFILLER_98_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7063_ _7063_/A _7161_/A vssd1 vssd1 vccd1 vccd1 _7064_/B sky130_fd_sc_hd__xnor2_1
XFILLER_98_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6014_ _5944_/Y _5916_/B _6169_/B vssd1 vssd1 vccd1 vccd1 _6014_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_100_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7965_ _7964_/A _7964_/B _7964_/C vssd1 vssd1 vccd1 vccd1 _7965_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_14_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7896_ _7831_/A _7831_/B _7895_/X vssd1 vssd1 vccd1 vccd1 _7982_/A sky130_fd_sc_hd__a21o_1
X_6916_ _6916_/A _7027_/A vssd1 vssd1 vccd1 vccd1 _6918_/B sky130_fd_sc_hd__xnor2_1
XFILLER_23_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6847_ _6976_/A _6976_/B _6846_/X vssd1 vssd1 vccd1 vccd1 _6892_/A sky130_fd_sc_hd__o21a_1
Xclkbuf_4_13_0_wb_clk_i clkbuf_3_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8785_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_50_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6778_ _6786_/A _6778_/B vssd1 vssd1 vccd1 vccd1 _6779_/B sky130_fd_sc_hd__xor2_1
X_8517_ _8453_/A _8517_/B vssd1 vssd1 vccd1 vccd1 _8518_/B sky130_fd_sc_hd__and2b_1
X_5729_ _5728_/B _5728_/C _5835_/A vssd1 vssd1 vccd1 vccd1 _5730_/C sky130_fd_sc_hd__o21ai_1
X_8448_ _8163_/A _7755_/X _8514_/B vssd1 vssd1 vccd1 vccd1 _8452_/A sky130_fd_sc_hd__a21o_1
X_8379_ _8514_/A _8514_/B vssd1 vssd1 vccd1 vccd1 _8461_/S sky130_fd_sc_hd__nor2_2
XFILLER_89_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8827__44 vssd1 vssd1 vccd1 vccd1 _8827__44/HI _8922_/A sky130_fd_sc_hd__conb_1
XFILLER_24_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7750_ _7913_/A _8172_/A vssd1 vssd1 vccd1 vccd1 _8450_/B sky130_fd_sc_hd__nor2_2
X_4962_ _5271_/B _4955_/X _4961_/X vssd1 vssd1 vccd1 vccd1 _4962_/X sky130_fd_sc_hd__o21a_1
X_7681_ _7681_/A _7681_/B vssd1 vssd1 vccd1 vccd1 _7693_/A sky130_fd_sc_hd__xnor2_2
X_4893_ _4921_/A _4912_/B vssd1 vssd1 vccd1 vccd1 _5283_/B sky130_fd_sc_hd__nor2_1
X_6701_ _6670_/A _6670_/B _6617_/A vssd1 vssd1 vccd1 vccd1 _6704_/A sky130_fd_sc_hd__a21o_1
X_6632_ _6632_/A _6632_/B vssd1 vssd1 vccd1 vccd1 _6774_/A sky130_fd_sc_hd__xnor2_2
X_6563_ _7587_/B _6563_/B vssd1 vssd1 vccd1 vccd1 _6568_/A sky130_fd_sc_hd__and2b_1
X_8302_ _8302_/A _8302_/B _8302_/C vssd1 vssd1 vccd1 vccd1 _8303_/B sky130_fd_sc_hd__nor3_1
X_5514_ _5552_/A _5526_/B vssd1 vssd1 vccd1 vccd1 _5853_/A sky130_fd_sc_hd__xnor2_4
X_6494_ _6497_/C _6494_/B vssd1 vssd1 vccd1 vccd1 _8734_/D sky130_fd_sc_hd__nor2_1
X_8233_ _8223_/A _8223_/B _8232_/X vssd1 vssd1 vccd1 vccd1 _8317_/A sky130_fd_sc_hd__a21boi_2
X_5445_ _5445_/A vssd1 vssd1 vccd1 vccd1 _5450_/A sky130_fd_sc_hd__clkbuf_2
X_8164_ _8270_/B _8066_/X _8064_/Y _8380_/A vssd1 vssd1 vccd1 vccd1 _8177_/A sky130_fd_sc_hd__a22o_1
X_7115_ _7157_/A _7157_/B vssd1 vssd1 vccd1 vccd1 _7530_/A sky130_fd_sc_hd__xor2_1
X_5376_ _6532_/D _5377_/C _5375_/Y vssd1 vssd1 vccd1 vccd1 _8692_/D sky130_fd_sc_hd__a21oi_1
XFILLER_87_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8095_ _8028_/A _8336_/A _8094_/Y vssd1 vssd1 vccd1 vccd1 _8096_/B sky130_fd_sc_hd__o21a_1
XFILLER_86_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7046_ _7370_/A vssd1 vssd1 vccd1 vccd1 _7484_/S sky130_fd_sc_hd__buf_2
XFILLER_74_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7948_ _7696_/A _8098_/A _8120_/A vssd1 vssd1 vccd1 vccd1 _7949_/B sky130_fd_sc_hd__a21oi_1
XFILLER_42_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7879_ _7904_/A _8182_/A vssd1 vssd1 vccd1 vccd1 _7880_/B sky130_fd_sc_hd__nor2_1
XFILLER_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5230_ _4960_/B _5226_/Y _5235_/A _5145_/Y _5229_/Y vssd1 vssd1 vccd1 vccd1 _5231_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5161_ _5136_/C _5158_/X _5159_/X _5033_/B _5259_/C vssd1 vssd1 vccd1 vccd1 _5170_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_96_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5092_ _5145_/B _5202_/A _5089_/X _5095_/C vssd1 vssd1 vccd1 vccd1 _5092_/X sky130_fd_sc_hd__a211o_1
X_8920_ _8920_/A _4405_/Y vssd1 vssd1 vccd1 vccd1 io_out[7] sky130_fd_sc_hd__ebufn_8
XFILLER_83_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7802_ _7818_/A _7802_/B vssd1 vssd1 vccd1 vccd1 _7897_/B sky130_fd_sc_hd__xnor2_1
X_8782_ _8785_/CLK _8782_/D vssd1 vssd1 vccd1 vccd1 _8782_/Q sky130_fd_sc_hd__dfxtp_1
X_5994_ _6085_/A _5994_/B vssd1 vssd1 vccd1 vccd1 _5995_/B sky130_fd_sc_hd__xnor2_1
XFILLER_37_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7733_ _7733_/A _7733_/B vssd1 vssd1 vccd1 vccd1 _7789_/B sky130_fd_sc_hd__nor2_4
XFILLER_24_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4945_ _4953_/C vssd1 vssd1 vccd1 vccd1 _4995_/C sky130_fd_sc_hd__clkbuf_2
X_7664_ _7775_/A _7644_/X _7663_/Y vssd1 vssd1 vccd1 vccd1 _8773_/D sky130_fd_sc_hd__a21o_1
X_4876_ _4902_/C _4879_/B vssd1 vssd1 vccd1 vccd1 _4889_/B sky130_fd_sc_hd__nand2_2
X_7595_ _8766_/Q vssd1 vssd1 vccd1 vccd1 _8612_/B sky130_fd_sc_hd__clkbuf_1
X_6615_ _8761_/Q _6615_/B vssd1 vssd1 vccd1 vccd1 _6617_/A sky130_fd_sc_hd__and2b_1
XFILLER_20_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6546_ _6541_/X _6543_/X _7583_/A _7585_/A vssd1 vssd1 vccd1 vccd1 _6546_/Y sky130_fd_sc_hd__a211oi_1
X_6477_ _6452_/A _6478_/C _6476_/Y vssd1 vssd1 vccd1 vccd1 _8729_/D sky130_fd_sc_hd__a21oi_1
X_8216_ _8214_/Y _8216_/B vssd1 vssd1 vccd1 vccd1 _8304_/B sky130_fd_sc_hd__and2b_1
X_5428_ _6427_/A _6420_/B _5423_/X _5427_/Y _4615_/A vssd1 vssd1 vccd1 vccd1 _5429_/A
+ sky130_fd_sc_hd__o311a_1
X_8147_ _8147_/A _8147_/B vssd1 vssd1 vccd1 vccd1 _8147_/Y sky130_fd_sc_hd__nand2_1
X_5359_ _8687_/Q _5359_/B vssd1 vssd1 vccd1 vccd1 _5365_/C sky130_fd_sc_hd__and2_1
X_8078_ _8078_/A _8078_/B vssd1 vssd1 vccd1 vccd1 _8079_/B sky130_fd_sc_hd__or2_1
XINSDIODE2_2 _5250_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7029_ _7301_/A _6813_/B _6933_/B _7028_/Y vssd1 vssd1 vccd1 vccd1 _7039_/A sky130_fd_sc_hd__a31o_1
XFILLER_74_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8788__5 vssd1 vssd1 vccd1 vccd1 _8788__5/HI _8883_/A sky130_fd_sc_hd__conb_1
XFILLER_99_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4730_ _4730_/A _5170_/A vssd1 vssd1 vccd1 vccd1 _4730_/Y sky130_fd_sc_hd__nand2_1
X_4661_ _8644_/Q _8645_/Q _4661_/C vssd1 vssd1 vccd1 vccd1 _4665_/B sky130_fd_sc_hd__and3_1
XFILLER_80_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6400_ _8574_/A _8717_/Q vssd1 vssd1 vccd1 vccd1 _6400_/Y sky130_fd_sc_hd__nor2_1
X_7380_ _7380_/A _7489_/B vssd1 vssd1 vccd1 vccd1 _7417_/B sky130_fd_sc_hd__xnor2_2
X_6331_ _6331_/A _6331_/B vssd1 vssd1 vccd1 vccd1 _6338_/A sky130_fd_sc_hd__xnor2_1
X_4592_ _4592_/A vssd1 vssd1 vccd1 vccd1 _8937_/A sky130_fd_sc_hd__clkbuf_2
X_6262_ _6262_/A _6262_/B vssd1 vssd1 vccd1 vccd1 _6263_/B sky130_fd_sc_hd__nand2_1
X_8001_ _8001_/A _8001_/B vssd1 vssd1 vccd1 vccd1 _8002_/C sky130_fd_sc_hd__xnor2_1
X_6193_ _6193_/A _6200_/A vssd1 vssd1 vccd1 vccd1 _6194_/B sky130_fd_sc_hd__xor2_1
X_5213_ _5271_/A _5204_/X _5212_/X _5130_/A vssd1 vssd1 vccd1 vccd1 _5213_/X sky130_fd_sc_hd__a211o_1
X_5144_ _5150_/A _5137_/X _5143_/Y _5271_/B vssd1 vssd1 vccd1 vccd1 _5144_/X sky130_fd_sc_hd__o211a_1
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5075_ _5163_/A vssd1 vssd1 vccd1 vccd1 _5221_/C sky130_fd_sc_hd__clkbuf_2
X_8903_ _8903_/A _4385_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[22] sky130_fd_sc_hd__ebufn_8
XFILLER_64_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5977_ _5977_/A _5977_/B vssd1 vssd1 vccd1 vccd1 _5977_/Y sky130_fd_sc_hd__nand2_1
XFILLER_12_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8765_ _8765_/CLK _8765_/D vssd1 vssd1 vccd1 vccd1 _8765_/Q sky130_fd_sc_hd__dfxtp_1
X_7716_ _7761_/A _7714_/B _7715_/X vssd1 vssd1 vccd1 vccd1 _7719_/A sky130_fd_sc_hd__a21bo_1
X_4928_ _5100_/B _5107_/B vssd1 vssd1 vccd1 vccd1 _5171_/B sky130_fd_sc_hd__and2_1
X_8696_ _8704_/CLK _8696_/D vssd1 vssd1 vccd1 vccd1 _8696_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7647_ _7652_/B _7648_/B vssd1 vssd1 vccd1 vccd1 _7647_/X sky130_fd_sc_hd__and2_1
XFILLER_60_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4859_ _4883_/A vssd1 vssd1 vccd1 vccd1 _4934_/A sky130_fd_sc_hd__clkbuf_2
X_7578_ _7585_/A _7578_/B vssd1 vssd1 vccd1 vccd1 _7578_/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6529_ _8699_/Q _8698_/Q _8703_/Q _8702_/Q vssd1 vssd1 vccd1 vccd1 _6529_/X sky130_fd_sc_hd__and4_1
XFILLER_69_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5900_ _6081_/A _5824_/B _5829_/B _5827_/X vssd1 vssd1 vccd1 vccd1 _6002_/A sky130_fd_sc_hd__a31oi_2
XFILLER_53_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6880_ _6894_/A _6894_/B vssd1 vssd1 vccd1 vccd1 _6889_/A sky130_fd_sc_hd__xnor2_1
XFILLER_46_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5831_ _5889_/A _5830_/B _5830_/C vssd1 vssd1 vccd1 vccd1 _5832_/C sky130_fd_sc_hd__a21o_1
XFILLER_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5762_ _5810_/A _5810_/B _5810_/C vssd1 vssd1 vccd1 vccd1 _5792_/A sky130_fd_sc_hd__nand3_1
X_8550_ _8550_/A _8550_/B vssd1 vssd1 vccd1 vccd1 _8550_/X sky130_fd_sc_hd__xor2_1
XFILLER_22_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4713_ _5283_/A vssd1 vssd1 vccd1 vccd1 _5042_/A sky130_fd_sc_hd__clkbuf_2
X_7501_ _7501_/A _7501_/B vssd1 vssd1 vccd1 vccd1 _7502_/B sky130_fd_sc_hd__xnor2_2
X_8481_ _8481_/A _8481_/B vssd1 vssd1 vccd1 vccd1 _8483_/B sky130_fd_sc_hd__xnor2_1
X_5693_ _5693_/A _5693_/B vssd1 vssd1 vccd1 vccd1 _5694_/B sky130_fd_sc_hd__and2_1
X_7432_ _7432_/A _7432_/B vssd1 vssd1 vccd1 vccd1 _7433_/B sky130_fd_sc_hd__xor2_4
XFILLER_30_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4644_ _8638_/Q _4643_/C _8639_/Q vssd1 vssd1 vccd1 vccd1 _4645_/C sky130_fd_sc_hd__a21o_1
X_4575_ _5305_/A vssd1 vssd1 vccd1 vccd1 _4584_/B sky130_fd_sc_hd__clkbuf_2
X_7363_ _7363_/A _7363_/B vssd1 vssd1 vccd1 vccd1 _7460_/S sky130_fd_sc_hd__nor2_2
X_6314_ _6314_/A _6314_/B vssd1 vssd1 vccd1 vccd1 _6315_/B sky130_fd_sc_hd__xnor2_1
X_7294_ _7294_/A _7294_/B vssd1 vssd1 vccd1 vccd1 _7294_/Y sky130_fd_sc_hd__nor2_1
X_6245_ _6243_/Y _6211_/B _6244_/Y vssd1 vssd1 vccd1 vccd1 _6300_/A sky130_fd_sc_hd__a21o_1
XFILLER_89_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6176_ _6252_/A _6246_/B vssd1 vssd1 vccd1 vccd1 _6177_/B sky130_fd_sc_hd__xnor2_1
XFILLER_69_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5127_ _5127_/A _5127_/B _5127_/C vssd1 vssd1 vccd1 vccd1 _5128_/B sky130_fd_sc_hd__or3_1
XFILLER_29_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5058_ _5190_/A _5281_/B vssd1 vssd1 vccd1 vccd1 _5059_/B sky130_fd_sc_hd__or2_1
XFILLER_29_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8748_ _8753_/CLK _8748_/D vssd1 vssd1 vccd1 vccd1 _8748_/Q sky130_fd_sc_hd__dfxtp_1
X_8679_ _8778_/CLK _8679_/D vssd1 vssd1 vccd1 vccd1 _8679_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4360_ _4363_/A vssd1 vssd1 vccd1 vccd1 _4360_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8872__89 vssd1 vssd1 vccd1 vccd1 _8872__89/HI _8981_/A sky130_fd_sc_hd__conb_1
X_6030_ _6053_/A _6030_/B vssd1 vssd1 vccd1 vccd1 _6045_/A sky130_fd_sc_hd__xnor2_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7981_ _7981_/A _7981_/B _7981_/C vssd1 vssd1 vccd1 vccd1 _7981_/X sky130_fd_sc_hd__and3_1
XFILLER_66_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6932_ _7028_/A _7028_/B vssd1 vssd1 vccd1 vccd1 _6933_/B sky130_fd_sc_hd__xor2_1
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6863_ _7020_/A _6863_/B _6863_/C vssd1 vssd1 vccd1 vccd1 _6876_/A sky130_fd_sc_hd__and3_1
X_5814_ _5744_/B _5744_/C _5744_/A vssd1 vssd1 vccd1 vccd1 _5832_/A sky130_fd_sc_hd__a21bo_1
X_8602_ _8602_/A _8602_/B vssd1 vssd1 vccd1 vccd1 _8603_/B sky130_fd_sc_hd__xor2_1
XFILLER_62_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6794_ _6910_/B vssd1 vssd1 vccd1 vccd1 _6863_/C sky130_fd_sc_hd__clkbuf_2
X_8533_ _8533_/A _8533_/B vssd1 vssd1 vccd1 vccd1 _8534_/B sky130_fd_sc_hd__xnor2_1
X_5745_ _5744_/A _5744_/B _5744_/C vssd1 vssd1 vccd1 vccd1 _5746_/C sky130_fd_sc_hd__a21o_1
X_8464_ _8279_/A _8393_/A _8512_/A vssd1 vssd1 vccd1 vccd1 _8465_/B sky130_fd_sc_hd__o21ba_1
X_5676_ _5676_/A _5676_/B vssd1 vssd1 vccd1 vccd1 _5677_/B sky130_fd_sc_hd__nand2_1
XFILLER_30_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4627_ _4640_/A vssd1 vssd1 vccd1 vccd1 _4672_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_7415_ _7415_/A _7491_/B vssd1 vssd1 vccd1 vccd1 _7419_/A sky130_fd_sc_hd__xnor2_1
X_8395_ _8394_/A _8394_/B _8394_/C vssd1 vssd1 vccd1 vccd1 _8396_/C sky130_fd_sc_hd__a21o_1
X_7346_ _7346_/A _7346_/B vssd1 vssd1 vccd1 vccd1 _7348_/C sky130_fd_sc_hd__xnor2_1
X_4558_ _4720_/A vssd1 vssd1 vccd1 vccd1 _4558_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_104_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7277_ _7276_/A _7276_/B _7276_/C vssd1 vssd1 vccd1 vccd1 _7278_/B sky130_fd_sc_hd__a21oi_1
X_4489_ _4489_/A vssd1 vssd1 vccd1 vccd1 _4489_/Y sky130_fd_sc_hd__inv_2
XFILLER_89_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6228_ _6228_/A vssd1 vssd1 vccd1 vccd1 _6228_/Y sky130_fd_sc_hd__inv_2
X_6159_ _6159_/A _6159_/B vssd1 vssd1 vccd1 vccd1 _6160_/B sky130_fd_sc_hd__xnor2_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5530_ _5530_/A _5530_/B vssd1 vssd1 vccd1 vccd1 _5682_/B sky130_fd_sc_hd__xor2_4
X_5461_ _5456_/B _5449_/X _5450_/X _5460_/Y vssd1 vssd1 vccd1 vccd1 _8709_/D sky130_fd_sc_hd__a22o_1
XFILLER_8_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4412_ _4413_/A vssd1 vssd1 vccd1 vccd1 _4412_/Y sky130_fd_sc_hd__inv_2
X_7200_ _7037_/A _7200_/B vssd1 vssd1 vccd1 vccd1 _7200_/X sky130_fd_sc_hd__and2b_1
X_8180_ _8180_/A _8246_/B vssd1 vssd1 vccd1 vccd1 _8187_/A sky130_fd_sc_hd__xnor2_4
X_5392_ _6567_/A vssd1 vssd1 vccd1 vccd1 _5392_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7131_ _7131_/A _7130_/A vssd1 vssd1 vccd1 vccd1 _7131_/X sky130_fd_sc_hd__or2b_1
XFILLER_59_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7062_ _7062_/A _7062_/B vssd1 vssd1 vccd1 vccd1 _7161_/A sky130_fd_sc_hd__xnor2_1
XFILLER_98_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6013_ _6171_/B vssd1 vssd1 vccd1 vccd1 _6228_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_100_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7964_ _7964_/A _7964_/B _7964_/C vssd1 vssd1 vccd1 vccd1 _7964_/X sky130_fd_sc_hd__and3_1
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6915_ _6870_/X _6875_/B _6871_/A vssd1 vssd1 vccd1 vccd1 _7027_/A sky130_fd_sc_hd__a21oi_2
X_7895_ _8450_/A _8568_/D _7895_/C vssd1 vssd1 vccd1 vccd1 _7895_/X sky130_fd_sc_hd__and3_1
XFILLER_35_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6846_ _6846_/A _6846_/B vssd1 vssd1 vccd1 vccd1 _6846_/X sky130_fd_sc_hd__or2_1
X_6777_ _6863_/B vssd1 vssd1 vccd1 vccd1 _6960_/B sky130_fd_sc_hd__clkbuf_2
X_8516_ _8452_/A _8516_/B vssd1 vssd1 vccd1 vccd1 _8518_/A sky130_fd_sc_hd__and2b_1
X_5728_ _5835_/A _5728_/B _5728_/C vssd1 vssd1 vccd1 vccd1 _5730_/B sky130_fd_sc_hd__or3_1
X_8447_ _8387_/B _8387_/C _8387_/A vssd1 vssd1 vccd1 vccd1 _8528_/A sky130_fd_sc_hd__a21bo_1
X_5659_ _5917_/A vssd1 vssd1 vccd1 vccd1 _6147_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_8378_ _8382_/A _8378_/B _8378_/C vssd1 vssd1 vccd1 vccd1 _8459_/B sky130_fd_sc_hd__or3_1
XFILLER_104_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7329_ _6682_/Y _7309_/B _7230_/B _7370_/B vssd1 vssd1 vccd1 vccd1 _7333_/A sky130_fd_sc_hd__a22o_1
XFILLER_89_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8842__59 vssd1 vssd1 vccd1 vccd1 _8842__59/HI _8951_/A sky130_fd_sc_hd__conb_1
XFILLER_76_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4961_ _5224_/B _5136_/B _5149_/C _4980_/C vssd1 vssd1 vccd1 vccd1 _4961_/X sky130_fd_sc_hd__or4_1
X_7680_ _7678_/X _7688_/A vssd1 vssd1 vccd1 vccd1 _7681_/B sky130_fd_sc_hd__and2b_1
X_6700_ _6825_/A _6949_/A vssd1 vssd1 vccd1 vccd1 _7105_/A sky130_fd_sc_hd__nor2_1
X_4892_ _4892_/A vssd1 vssd1 vccd1 vccd1 _4912_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_32_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6631_ _6645_/A _6647_/B _6630_/X vssd1 vssd1 vccd1 vccd1 _6632_/B sky130_fd_sc_hd__a21o_2
X_8301_ _8302_/A _8302_/B _8302_/C vssd1 vssd1 vccd1 vccd1 _8303_/A sky130_fd_sc_hd__o21a_1
X_6562_ _6562_/A vssd1 vssd1 vccd1 vccd1 _7587_/B sky130_fd_sc_hd__clkbuf_2
X_5513_ _5698_/A vssd1 vssd1 vccd1 vccd1 _5852_/A sky130_fd_sc_hd__clkbuf_2
X_6493_ _8734_/Q _6491_/A _6465_/X vssd1 vssd1 vccd1 vccd1 _6494_/B sky130_fd_sc_hd__o21ai_1
X_8232_ _8232_/A _8207_/B vssd1 vssd1 vccd1 vccd1 _8232_/X sky130_fd_sc_hd__or2b_1
X_5444_ _6563_/B _5462_/A _5462_/B vssd1 vssd1 vccd1 vccd1 _5445_/A sky130_fd_sc_hd__and3_1
X_8163_ _8163_/A _8163_/B vssd1 vssd1 vccd1 vccd1 _8272_/C sky130_fd_sc_hd__nor2_1
X_7114_ _7111_/A _7111_/B _7113_/X vssd1 vssd1 vccd1 vccd1 _7157_/B sky130_fd_sc_hd__a21oi_1
X_5375_ _6532_/D _5377_/C _5409_/A vssd1 vssd1 vccd1 vccd1 _5375_/Y sky130_fd_sc_hd__o21ai_1
X_8094_ _8239_/A _8420_/A vssd1 vssd1 vccd1 vccd1 _8094_/Y sky130_fd_sc_hd__nand2_1
XFILLER_59_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7045_ _7469_/A _7228_/B vssd1 vssd1 vccd1 vccd1 _7370_/A sky130_fd_sc_hd__xnor2_1
XFILLER_86_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7947_ _7845_/A _7845_/B _8120_/A _7696_/A vssd1 vssd1 vccd1 vccd1 _8044_/A sky130_fd_sc_hd__o211a_2
XFILLER_70_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7878_ _7940_/A _8103_/A _7878_/C vssd1 vssd1 vccd1 vccd1 _8567_/A sky130_fd_sc_hd__and3_1
X_6829_ _6829_/A _6829_/B vssd1 vssd1 vccd1 vccd1 _6973_/B sky130_fd_sc_hd__xnor2_2
XFILLER_12_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5160_ _5160_/A vssd1 vssd1 vccd1 vccd1 _5259_/C sky130_fd_sc_hd__clkbuf_2
X_5091_ _5138_/A _5120_/B _5099_/D vssd1 vssd1 vccd1 vccd1 _5095_/C sky130_fd_sc_hd__or3_1
XFILLER_37_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7801_ _8273_/A _8165_/C _7768_/A _7800_/Y vssd1 vssd1 vccd1 vccd1 _7802_/B sky130_fd_sc_hd__o211a_1
X_8781_ _8783_/CLK _8781_/D vssd1 vssd1 vccd1 vccd1 _8781_/Q sky130_fd_sc_hd__dfxtp_1
X_5993_ _5993_/A _5993_/B vssd1 vssd1 vccd1 vccd1 _6085_/A sky130_fd_sc_hd__or2_2
XFILLER_52_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7732_ _8658_/Q _8782_/Q vssd1 vssd1 vccd1 vccd1 _7733_/B sky130_fd_sc_hd__and2b_1
XFILLER_52_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4944_ _4957_/A _4966_/A vssd1 vssd1 vccd1 vccd1 _4953_/C sky130_fd_sc_hd__or2_1
X_7663_ _7644_/X _7662_/Y _7624_/X vssd1 vssd1 vccd1 vccd1 _7663_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_32_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4875_ _5298_/B _5298_/C vssd1 vssd1 vccd1 vccd1 _4879_/B sky130_fd_sc_hd__nor2_1
X_7594_ _8782_/Q vssd1 vssd1 vccd1 vccd1 _8605_/A sky130_fd_sc_hd__inv_2
X_6614_ _6648_/A _6637_/B _6613_/X vssd1 vssd1 vccd1 vccd1 _6670_/A sky130_fd_sc_hd__a21o_4
XFILLER_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6545_ _8763_/Q vssd1 vssd1 vccd1 vccd1 _7585_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_8215_ _8214_/A _8214_/C _8214_/B vssd1 vssd1 vccd1 vccd1 _8216_/B sky130_fd_sc_hd__o21ai_1
X_6476_ _6452_/A _6478_/C _6524_/B vssd1 vssd1 vccd1 vccd1 _6476_/Y sky130_fd_sc_hd__o21ai_1
X_5427_ _6433_/A _5440_/C _6427_/B vssd1 vssd1 vccd1 vccd1 _5427_/Y sky130_fd_sc_hd__o21ai_1
X_8146_ _8133_/A _8133_/B _8145_/X vssd1 vssd1 vccd1 vccd1 _8229_/A sky130_fd_sc_hd__a21oi_2
XFILLER_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5358_ _5358_/A vssd1 vssd1 vccd1 vccd1 _8686_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8077_ _8078_/A _8078_/B vssd1 vssd1 vccd1 vccd1 _8185_/B sky130_fd_sc_hd__nand2_1
XFILLER_58_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_3 _5128_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7028_ _7028_/A _7028_/B vssd1 vssd1 vccd1 vccd1 _7028_/Y sky130_fd_sc_hd__nor2_1
X_5289_ _4964_/X _5087_/B _5188_/D _5288_/X vssd1 vssd1 vccd1 vccd1 _5289_/X sky130_fd_sc_hd__o31a_1
XFILLER_74_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8979_ _8979_/A _4474_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[28] sky130_fd_sc_hd__ebufn_8
XFILLER_82_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8812__29 vssd1 vssd1 vccd1 vccd1 _8812__29/HI _8907_/A sky130_fd_sc_hd__conb_1
XFILLER_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4660_ _8644_/Q _4661_/C _4659_/Y vssd1 vssd1 vccd1 vccd1 _8644_/D sky130_fd_sc_hd__a21oi_1
XFILLER_80_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6330_ _6330_/A _6330_/B vssd1 vssd1 vccd1 vccd1 _6331_/B sky130_fd_sc_hd__xnor2_2
X_4591_ _8683_/Q _4595_/B vssd1 vssd1 vccd1 vccd1 _4592_/A sky130_fd_sc_hd__and2_1
X_6261_ _6262_/A _5595_/Y _6264_/A vssd1 vssd1 vccd1 vccd1 _6265_/A sky130_fd_sc_hd__a21o_1
X_8000_ _8261_/A _7925_/A _7999_/X vssd1 vssd1 vccd1 vccd1 _8001_/B sky130_fd_sc_hd__a21oi_1
X_6192_ _6192_/A _6192_/B vssd1 vssd1 vccd1 vccd1 _6200_/A sky130_fd_sc_hd__nor2_1
X_5212_ _4965_/X _5205_/X _5211_/X _5136_/C _4558_/X vssd1 vssd1 vccd1 vccd1 _5212_/X
+ sky130_fd_sc_hd__o221a_1
X_5143_ _5140_/Y _5141_/X _5142_/Y vssd1 vssd1 vccd1 vccd1 _5143_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_84_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5074_ _5277_/B _5074_/B _5141_/C vssd1 vssd1 vccd1 vccd1 _5227_/A sky130_fd_sc_hd__or3b_2
X_8902_ _8902_/A _4384_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[21] sky130_fd_sc_hd__ebufn_8
XFILLER_71_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5976_ _5905_/A _5905_/B _5975_/Y vssd1 vssd1 vccd1 vccd1 _6001_/A sky130_fd_sc_hd__o21a_1
XFILLER_25_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8764_ _8784_/CLK _8764_/D vssd1 vssd1 vccd1 vccd1 _8764_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7715_ _7764_/A _7764_/B vssd1 vssd1 vccd1 vccd1 _7715_/X sky130_fd_sc_hd__or2_1
XFILLER_52_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8695_ _8704_/CLK _8695_/D vssd1 vssd1 vccd1 vccd1 _8695_/Q sky130_fd_sc_hd__dfxtp_1
X_4927_ _4927_/A _4927_/B _5298_/C vssd1 vssd1 vccd1 vccd1 _5107_/B sky130_fd_sc_hd__and3_1
X_7646_ _7638_/A _7640_/B _7638_/B vssd1 vssd1 vccd1 vccd1 _7648_/B sky130_fd_sc_hd__o21ba_1
X_4858_ _7684_/B _5501_/B _4927_/A vssd1 vssd1 vccd1 vccd1 _4883_/A sky130_fd_sc_hd__or3_1
X_7577_ _6569_/A _7586_/S _7575_/X _7576_/X vssd1 vssd1 vccd1 vccd1 _8763_/D sky130_fd_sc_hd__a31o_1
X_4789_ _4791_/A vssd1 vssd1 vccd1 vccd1 _5334_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_8878__95 vssd1 vssd1 vccd1 vccd1 _8878__95/HI _8987_/A sky130_fd_sc_hd__conb_1
X_6528_ _8691_/Q _8690_/Q _6528_/C _8694_/Q vssd1 vssd1 vccd1 vccd1 _6535_/B sky130_fd_sc_hd__nand4_1
XFILLER_69_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6459_ _7622_/A _7622_/B vssd1 vssd1 vccd1 vccd1 _8628_/A sky130_fd_sc_hd__or2_2
XFILLER_0_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8129_ _8222_/A _8129_/B vssd1 vssd1 vccd1 vccd1 _8131_/B sky130_fd_sc_hd__nand2_1
XFILLER_102_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8790__7 vssd1 vssd1 vccd1 vccd1 _8790__7/HI _8885_/A sky130_fd_sc_hd__conb_1
XFILLER_18_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5830_ _5889_/A _5830_/B _5830_/C vssd1 vssd1 vccd1 vccd1 _5889_/B sky130_fd_sc_hd__nand3_1
X_5761_ _6071_/A _6197_/A _5760_/C _5760_/D vssd1 vssd1 vccd1 vccd1 _5810_/C sky130_fd_sc_hd__a22o_1
XFILLER_61_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8480_ _8480_/A _8480_/B vssd1 vssd1 vccd1 vccd1 _8483_/A sky130_fd_sc_hd__or2_1
X_7500_ _7500_/A _7500_/B vssd1 vssd1 vccd1 vccd1 _7501_/B sky130_fd_sc_hd__xnor2_1
X_4712_ _8652_/Q vssd1 vssd1 vccd1 vccd1 _5283_/A sky130_fd_sc_hd__inv_2
X_5692_ _5693_/A _5693_/B vssd1 vssd1 vccd1 vccd1 _5694_/A sky130_fd_sc_hd__nor2_1
X_7431_ _7442_/A _7442_/B vssd1 vssd1 vccd1 vccd1 _7432_/B sky130_fd_sc_hd__xor2_4
XFILLER_30_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4643_ _8638_/Q _8639_/Q _4643_/C vssd1 vssd1 vccd1 vccd1 _4647_/B sky130_fd_sc_hd__and3_1
X_7362_ _7333_/A _7360_/Y _7361_/X vssd1 vssd1 vccd1 vccd1 _7462_/A sky130_fd_sc_hd__a21bo_1
X_4574_ _4574_/A _4574_/B _4574_/C _4574_/D vssd1 vssd1 vccd1 vccd1 _5305_/A sky130_fd_sc_hd__and4_1
X_6313_ _6313_/A _6313_/B vssd1 vssd1 vccd1 vccd1 _6314_/B sky130_fd_sc_hd__xnor2_1
X_7293_ _7293_/A _7293_/B vssd1 vssd1 vccd1 vccd1 _7427_/A sky130_fd_sc_hd__xor2_2
X_6244_ _6244_/A _6244_/B vssd1 vssd1 vccd1 vccd1 _6244_/Y sky130_fd_sc_hd__nor2_1
XFILLER_103_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6175_ _6175_/A _6175_/B vssd1 vssd1 vccd1 vccd1 _6246_/B sky130_fd_sc_hd__xnor2_1
XFILLER_69_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5126_ _8654_/Q _5138_/A _5159_/D _5126_/D vssd1 vssd1 vccd1 vccd1 _5127_/C sky130_fd_sc_hd__or4_1
XFILLER_57_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5057_ _5209_/A vssd1 vssd1 vccd1 vccd1 _5250_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_53_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5959_ _5959_/A _5962_/B vssd1 vssd1 vccd1 vccd1 _5965_/A sky130_fd_sc_hd__or2_1
XFILLER_52_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8747_ _8753_/CLK _8747_/D vssd1 vssd1 vccd1 vccd1 _8747_/Q sky130_fd_sc_hd__dfxtp_1
X_8678_ _8778_/CLK _8678_/D vssd1 vssd1 vccd1 vccd1 _8678_/Q sky130_fd_sc_hd__dfxtp_1
X_7629_ _8768_/Q vssd1 vssd1 vccd1 vccd1 _7672_/A sky130_fd_sc_hd__inv_2
XFILLER_20_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7980_ _7887_/Y _8582_/A _7979_/X vssd1 vssd1 vccd1 vccd1 _8578_/A sky130_fd_sc_hd__a21oi_1
XFILLER_54_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6931_ _6943_/A _7303_/A vssd1 vssd1 vccd1 vccd1 _7028_/B sky130_fd_sc_hd__xnor2_1
XFILLER_62_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6862_ _6765_/A _6866_/C _7400_/B _6863_/C vssd1 vssd1 vccd1 vccd1 _6862_/X sky130_fd_sc_hd__a22o_1
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5813_ _5756_/B _5756_/C _5756_/A vssd1 vssd1 vccd1 vccd1 _5843_/A sky130_fd_sc_hd__a21bo_1
XFILLER_62_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8601_ _7739_/A _8595_/B _8594_/A vssd1 vssd1 vccd1 vccd1 _8602_/B sky130_fd_sc_hd__o21ai_1
XFILLER_22_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8532_ _8532_/A _8532_/B vssd1 vssd1 vccd1 vccd1 _8533_/B sky130_fd_sc_hd__xnor2_1
X_6793_ _6793_/A _7262_/B _6793_/C vssd1 vssd1 vccd1 vccd1 _6804_/A sky130_fd_sc_hd__or3_1
X_5744_ _5744_/A _5744_/B _5744_/C vssd1 vssd1 vccd1 vccd1 _5746_/B sky130_fd_sc_hd__nand3_1
X_8463_ _8463_/A _8463_/B _8463_/C vssd1 vssd1 vccd1 vccd1 _8512_/A sky130_fd_sc_hd__and3_1
X_5675_ _5715_/A _5674_/C _5679_/A vssd1 vssd1 vccd1 vccd1 _5676_/B sky130_fd_sc_hd__o21ai_1
X_8394_ _8394_/A _8394_/B _8394_/C vssd1 vssd1 vccd1 vccd1 _8396_/B sky130_fd_sc_hd__nand3_1
X_7414_ _7123_/B _7501_/A _7281_/A _7413_/Y vssd1 vssd1 vccd1 vccd1 _7491_/B sky130_fd_sc_hd__a22o_1
X_4626_ _8634_/Q _4631_/C vssd1 vssd1 vccd1 vccd1 _4630_/A sky130_fd_sc_hd__and2_1
X_8848__65 vssd1 vssd1 vccd1 vccd1 _8848__65/HI _8957_/A sky130_fd_sc_hd__conb_1
X_7345_ _7345_/A _7345_/B vssd1 vssd1 vccd1 vccd1 _7346_/B sky130_fd_sc_hd__xor2_1
X_4557_ _4733_/C vssd1 vssd1 vccd1 vccd1 _4720_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_103_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4488_ _4489_/A vssd1 vssd1 vccd1 vccd1 _4488_/Y sky130_fd_sc_hd__inv_2
XFILLER_89_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7276_ _7276_/A _7276_/B _7276_/C vssd1 vssd1 vccd1 vccd1 _7278_/A sky130_fd_sc_hd__and3_1
XFILLER_89_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6227_ _6227_/A _6227_/B vssd1 vssd1 vccd1 vccd1 _6232_/A sky130_fd_sc_hd__nand2_1
X_6158_ _6158_/A _6158_/B vssd1 vssd1 vccd1 vccd1 _6159_/B sky130_fd_sc_hd__nand2_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5109_ _5117_/B _5141_/D vssd1 vssd1 vccd1 vccd1 _5197_/A sky130_fd_sc_hd__nand2_1
X_6089_ _6089_/A vssd1 vssd1 vccd1 vccd1 _6278_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_72_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5460_ _5460_/A _5460_/B vssd1 vssd1 vccd1 vccd1 _5460_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_8_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4411_ _4413_/A vssd1 vssd1 vccd1 vccd1 _4411_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5391_ _8697_/Q _5395_/C vssd1 vssd1 vccd1 vccd1 _5394_/A sky130_fd_sc_hd__and2_1
X_7130_ _7130_/A _7131_/A vssd1 vssd1 vccd1 vccd1 _7137_/B sky130_fd_sc_hd__xor2_1
X_7061_ _7061_/A _7061_/B vssd1 vssd1 vccd1 vccd1 _7062_/B sky130_fd_sc_hd__xor2_1
X_6012_ _6012_/A _6165_/B vssd1 vssd1 vccd1 vccd1 _6171_/B sky130_fd_sc_hd__or2_1
.ends

