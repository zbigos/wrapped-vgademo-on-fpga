magic
tech sky130A
magscale 1 2
timestamp 1647765932
<< obsli1 >>
rect 1104 527 58880 57681
<< obsm1 >>
rect 566 416 59326 57712
<< metal2 >>
rect 542 59200 654 60000
rect 1738 59200 1850 60000
rect 2934 59200 3046 60000
rect 4130 59200 4242 60000
rect 5418 59200 5530 60000
rect 6614 59200 6726 60000
rect 7810 59200 7922 60000
rect 9098 59200 9210 60000
rect 10294 59200 10406 60000
rect 11490 59200 11602 60000
rect 12778 59200 12890 60000
rect 13974 59200 14086 60000
rect 15170 59200 15282 60000
rect 16366 59200 16478 60000
rect 17654 59200 17766 60000
rect 18850 59200 18962 60000
rect 20046 59200 20158 60000
rect 21334 59200 21446 60000
rect 22530 59200 22642 60000
rect 23726 59200 23838 60000
rect 25014 59200 25126 60000
rect 26210 59200 26322 60000
rect 27406 59200 27518 60000
rect 28694 59200 28806 60000
rect 29890 59200 30002 60000
rect 31086 59200 31198 60000
rect 32282 59200 32394 60000
rect 33570 59200 33682 60000
rect 34766 59200 34878 60000
rect 35962 59200 36074 60000
rect 37250 59200 37362 60000
rect 38446 59200 38558 60000
rect 39642 59200 39754 60000
rect 40930 59200 41042 60000
rect 42126 59200 42238 60000
rect 43322 59200 43434 60000
rect 44610 59200 44722 60000
rect 45806 59200 45918 60000
rect 47002 59200 47114 60000
rect 48198 59200 48310 60000
rect 49486 59200 49598 60000
rect 50682 59200 50794 60000
rect 51878 59200 51990 60000
rect 53166 59200 53278 60000
rect 54362 59200 54474 60000
rect 55558 59200 55670 60000
rect 56846 59200 56958 60000
rect 58042 59200 58154 60000
rect 59238 59200 59350 60000
rect 2658 0 2770 800
rect 8086 0 8198 800
rect 13514 0 13626 800
rect 18942 0 19054 800
rect 24462 0 24574 800
rect 29890 0 30002 800
rect 35318 0 35430 800
rect 40746 0 40858 800
rect 46266 0 46378 800
rect 51694 0 51806 800
rect 57122 0 57234 800
<< obsm2 >>
rect 710 59144 1682 59537
rect 1906 59144 2878 59537
rect 3102 59144 4074 59537
rect 4298 59144 5362 59537
rect 5586 59144 6558 59537
rect 6782 59144 7754 59537
rect 7978 59144 9042 59537
rect 9266 59144 10238 59537
rect 10462 59144 11434 59537
rect 11658 59144 12722 59537
rect 12946 59144 13918 59537
rect 14142 59144 15114 59537
rect 15338 59144 16310 59537
rect 16534 59144 17598 59537
rect 17822 59144 18794 59537
rect 19018 59144 19990 59537
rect 20214 59144 21278 59537
rect 21502 59144 22474 59537
rect 22698 59144 23670 59537
rect 23894 59144 24958 59537
rect 25182 59144 26154 59537
rect 26378 59144 27350 59537
rect 27574 59144 28638 59537
rect 28862 59144 29834 59537
rect 30058 59144 31030 59537
rect 31254 59144 32226 59537
rect 32450 59144 33514 59537
rect 33738 59144 34710 59537
rect 34934 59144 35906 59537
rect 36130 59144 37194 59537
rect 37418 59144 38390 59537
rect 38614 59144 39586 59537
rect 39810 59144 40874 59537
rect 41098 59144 42070 59537
rect 42294 59144 43266 59537
rect 43490 59144 44554 59537
rect 44778 59144 45750 59537
rect 45974 59144 46946 59537
rect 47170 59144 48142 59537
rect 48366 59144 49430 59537
rect 49654 59144 50626 59537
rect 50850 59144 51822 59537
rect 52046 59144 53110 59537
rect 53334 59144 54306 59537
rect 54530 59144 55502 59537
rect 55726 59144 56790 59537
rect 57014 59144 57986 59537
rect 58210 59144 59182 59537
rect 572 856 59320 59144
rect 572 410 2602 856
rect 2826 410 8030 856
rect 8254 410 13458 856
rect 13682 410 18886 856
rect 19110 410 24406 856
rect 24630 410 29834 856
rect 30058 410 35262 856
rect 35486 410 40690 856
rect 40914 410 46210 856
rect 46434 410 51638 856
rect 51862 410 57066 856
rect 57290 410 59320 856
<< metal3 >>
rect 0 59380 800 59620
rect 59200 59380 60000 59620
rect 0 58564 800 58804
rect 59200 58564 60000 58804
rect 0 57748 800 57988
rect 59200 57884 60000 58124
rect 0 56932 800 57172
rect 59200 57068 60000 57308
rect 0 56116 800 56356
rect 59200 56388 60000 56628
rect 0 55300 800 55540
rect 59200 55572 60000 55812
rect 0 54484 800 54724
rect 59200 54756 60000 54996
rect 59200 54076 60000 54316
rect 0 53668 800 53908
rect 59200 53260 60000 53500
rect 0 52852 800 53092
rect 59200 52580 60000 52820
rect 0 52036 800 52276
rect 59200 51764 60000 52004
rect 0 51220 800 51460
rect 59200 51084 60000 51324
rect 0 50404 800 50644
rect 59200 50268 60000 50508
rect 0 49588 800 49828
rect 59200 49452 60000 49692
rect 0 48772 800 49012
rect 59200 48772 60000 49012
rect 0 47956 800 48196
rect 59200 47956 60000 48196
rect 0 47140 800 47380
rect 59200 47276 60000 47516
rect 0 46324 800 46564
rect 59200 46460 60000 46700
rect 0 45508 800 45748
rect 59200 45644 60000 45884
rect 0 44692 800 44932
rect 59200 44964 60000 45204
rect 0 43876 800 44116
rect 59200 44148 60000 44388
rect 59200 43468 60000 43708
rect 0 43060 800 43300
rect 59200 42652 60000 42892
rect 0 42244 800 42484
rect 59200 41972 60000 42212
rect 0 41428 800 41668
rect 59200 41156 60000 41396
rect 0 40612 800 40852
rect 59200 40340 60000 40580
rect 0 39660 800 39900
rect 59200 39660 60000 39900
rect 0 38844 800 39084
rect 59200 38844 60000 39084
rect 0 38028 800 38268
rect 59200 38164 60000 38404
rect 0 37212 800 37452
rect 59200 37348 60000 37588
rect 0 36396 800 36636
rect 59200 36532 60000 36772
rect 0 35580 800 35820
rect 59200 35852 60000 36092
rect 0 34764 800 35004
rect 59200 35036 60000 35276
rect 59200 34356 60000 34596
rect 0 33948 800 34188
rect 59200 33540 60000 33780
rect 0 33132 800 33372
rect 59200 32860 60000 33100
rect 0 32316 800 32556
rect 59200 32044 60000 32284
rect 0 31500 800 31740
rect 59200 31228 60000 31468
rect 0 30684 800 30924
rect 59200 30548 60000 30788
rect 0 29868 800 30108
rect 59200 29732 60000 29972
rect 0 29052 800 29292
rect 59200 29052 60000 29292
rect 0 28236 800 28476
rect 59200 28236 60000 28476
rect 0 27420 800 27660
rect 59200 27420 60000 27660
rect 0 26604 800 26844
rect 59200 26740 60000 26980
rect 0 25788 800 26028
rect 59200 25924 60000 26164
rect 0 24972 800 25212
rect 59200 25244 60000 25484
rect 0 24156 800 24396
rect 59200 24428 60000 24668
rect 59200 23748 60000 23988
rect 0 23340 800 23580
rect 59200 22932 60000 23172
rect 0 22524 800 22764
rect 59200 22116 60000 22356
rect 0 21708 800 21948
rect 59200 21436 60000 21676
rect 0 20892 800 21132
rect 59200 20620 60000 20860
rect 0 19940 800 20180
rect 59200 19940 60000 20180
rect 0 19124 800 19364
rect 59200 19124 60000 19364
rect 0 18308 800 18548
rect 59200 18308 60000 18548
rect 0 17492 800 17732
rect 59200 17628 60000 17868
rect 0 16676 800 16916
rect 59200 16812 60000 17052
rect 0 15860 800 16100
rect 59200 16132 60000 16372
rect 0 15044 800 15284
rect 59200 15316 60000 15556
rect 59200 14636 60000 14876
rect 0 14228 800 14468
rect 59200 13820 60000 14060
rect 0 13412 800 13652
rect 59200 13004 60000 13244
rect 0 12596 800 12836
rect 59200 12324 60000 12564
rect 0 11780 800 12020
rect 59200 11508 60000 11748
rect 0 10964 800 11204
rect 59200 10828 60000 11068
rect 0 10148 800 10388
rect 59200 10012 60000 10252
rect 0 9332 800 9572
rect 59200 9196 60000 9436
rect 0 8516 800 8756
rect 59200 8516 60000 8756
rect 0 7700 800 7940
rect 59200 7700 60000 7940
rect 0 6884 800 7124
rect 59200 7020 60000 7260
rect 0 6068 800 6308
rect 59200 6204 60000 6444
rect 0 5252 800 5492
rect 59200 5524 60000 5764
rect 0 4436 800 4676
rect 59200 4708 60000 4948
rect 0 3620 800 3860
rect 59200 3892 60000 4132
rect 59200 3212 60000 3452
rect 0 2804 800 3044
rect 59200 2396 60000 2636
rect 0 1988 800 2228
rect 59200 1716 60000 1956
rect 0 1172 800 1412
rect 59200 900 60000 1140
rect 0 356 800 596
rect 59200 220 60000 460
<< obsm3 >>
rect 880 59300 59120 59533
rect 800 58884 59200 59300
rect 880 58484 59120 58884
rect 800 58204 59200 58484
rect 800 58068 59120 58204
rect 880 57804 59120 58068
rect 880 57668 59200 57804
rect 800 57388 59200 57668
rect 800 57252 59120 57388
rect 880 56988 59120 57252
rect 880 56852 59200 56988
rect 800 56708 59200 56852
rect 800 56436 59120 56708
rect 880 56308 59120 56436
rect 880 56036 59200 56308
rect 800 55892 59200 56036
rect 800 55620 59120 55892
rect 880 55492 59120 55620
rect 880 55220 59200 55492
rect 800 55076 59200 55220
rect 800 54804 59120 55076
rect 880 54676 59120 54804
rect 880 54404 59200 54676
rect 800 54396 59200 54404
rect 800 53996 59120 54396
rect 800 53988 59200 53996
rect 880 53588 59200 53988
rect 800 53580 59200 53588
rect 800 53180 59120 53580
rect 800 53172 59200 53180
rect 880 52900 59200 53172
rect 880 52772 59120 52900
rect 800 52500 59120 52772
rect 800 52356 59200 52500
rect 880 52084 59200 52356
rect 880 51956 59120 52084
rect 800 51684 59120 51956
rect 800 51540 59200 51684
rect 880 51404 59200 51540
rect 880 51140 59120 51404
rect 800 51004 59120 51140
rect 800 50724 59200 51004
rect 880 50588 59200 50724
rect 880 50324 59120 50588
rect 800 50188 59120 50324
rect 800 49908 59200 50188
rect 880 49772 59200 49908
rect 880 49508 59120 49772
rect 800 49372 59120 49508
rect 800 49092 59200 49372
rect 880 48692 59120 49092
rect 800 48276 59200 48692
rect 880 47876 59120 48276
rect 800 47596 59200 47876
rect 800 47460 59120 47596
rect 880 47196 59120 47460
rect 880 47060 59200 47196
rect 800 46780 59200 47060
rect 800 46644 59120 46780
rect 880 46380 59120 46644
rect 880 46244 59200 46380
rect 800 45964 59200 46244
rect 800 45828 59120 45964
rect 880 45564 59120 45828
rect 880 45428 59200 45564
rect 800 45284 59200 45428
rect 800 45012 59120 45284
rect 880 44884 59120 45012
rect 880 44612 59200 44884
rect 800 44468 59200 44612
rect 800 44196 59120 44468
rect 880 44068 59120 44196
rect 880 43796 59200 44068
rect 800 43788 59200 43796
rect 800 43388 59120 43788
rect 800 43380 59200 43388
rect 880 42980 59200 43380
rect 800 42972 59200 42980
rect 800 42572 59120 42972
rect 800 42564 59200 42572
rect 880 42292 59200 42564
rect 880 42164 59120 42292
rect 800 41892 59120 42164
rect 800 41748 59200 41892
rect 880 41476 59200 41748
rect 880 41348 59120 41476
rect 800 41076 59120 41348
rect 800 40932 59200 41076
rect 880 40660 59200 40932
rect 880 40532 59120 40660
rect 800 40260 59120 40532
rect 800 39980 59200 40260
rect 880 39580 59120 39980
rect 800 39164 59200 39580
rect 880 38764 59120 39164
rect 800 38484 59200 38764
rect 800 38348 59120 38484
rect 880 38084 59120 38348
rect 880 37948 59200 38084
rect 800 37668 59200 37948
rect 800 37532 59120 37668
rect 880 37268 59120 37532
rect 880 37132 59200 37268
rect 800 36852 59200 37132
rect 800 36716 59120 36852
rect 880 36452 59120 36716
rect 880 36316 59200 36452
rect 800 36172 59200 36316
rect 800 35900 59120 36172
rect 880 35772 59120 35900
rect 880 35500 59200 35772
rect 800 35356 59200 35500
rect 800 35084 59120 35356
rect 880 34956 59120 35084
rect 880 34684 59200 34956
rect 800 34676 59200 34684
rect 800 34276 59120 34676
rect 800 34268 59200 34276
rect 880 33868 59200 34268
rect 800 33860 59200 33868
rect 800 33460 59120 33860
rect 800 33452 59200 33460
rect 880 33180 59200 33452
rect 880 33052 59120 33180
rect 800 32780 59120 33052
rect 800 32636 59200 32780
rect 880 32364 59200 32636
rect 880 32236 59120 32364
rect 800 31964 59120 32236
rect 800 31820 59200 31964
rect 880 31548 59200 31820
rect 880 31420 59120 31548
rect 800 31148 59120 31420
rect 800 31004 59200 31148
rect 880 30868 59200 31004
rect 880 30604 59120 30868
rect 800 30468 59120 30604
rect 800 30188 59200 30468
rect 880 30052 59200 30188
rect 880 29788 59120 30052
rect 800 29652 59120 29788
rect 800 29372 59200 29652
rect 880 28972 59120 29372
rect 800 28556 59200 28972
rect 880 28156 59120 28556
rect 800 27740 59200 28156
rect 880 27340 59120 27740
rect 800 27060 59200 27340
rect 800 26924 59120 27060
rect 880 26660 59120 26924
rect 880 26524 59200 26660
rect 800 26244 59200 26524
rect 800 26108 59120 26244
rect 880 25844 59120 26108
rect 880 25708 59200 25844
rect 800 25564 59200 25708
rect 800 25292 59120 25564
rect 880 25164 59120 25292
rect 880 24892 59200 25164
rect 800 24748 59200 24892
rect 800 24476 59120 24748
rect 880 24348 59120 24476
rect 880 24076 59200 24348
rect 800 24068 59200 24076
rect 800 23668 59120 24068
rect 800 23660 59200 23668
rect 880 23260 59200 23660
rect 800 23252 59200 23260
rect 800 22852 59120 23252
rect 800 22844 59200 22852
rect 880 22444 59200 22844
rect 800 22436 59200 22444
rect 800 22036 59120 22436
rect 800 22028 59200 22036
rect 880 21756 59200 22028
rect 880 21628 59120 21756
rect 800 21356 59120 21628
rect 800 21212 59200 21356
rect 880 20940 59200 21212
rect 880 20812 59120 20940
rect 800 20540 59120 20812
rect 800 20260 59200 20540
rect 880 19860 59120 20260
rect 800 19444 59200 19860
rect 880 19044 59120 19444
rect 800 18628 59200 19044
rect 880 18228 59120 18628
rect 800 17948 59200 18228
rect 800 17812 59120 17948
rect 880 17548 59120 17812
rect 880 17412 59200 17548
rect 800 17132 59200 17412
rect 800 16996 59120 17132
rect 880 16732 59120 16996
rect 880 16596 59200 16732
rect 800 16452 59200 16596
rect 800 16180 59120 16452
rect 880 16052 59120 16180
rect 880 15780 59200 16052
rect 800 15636 59200 15780
rect 800 15364 59120 15636
rect 880 15236 59120 15364
rect 880 14964 59200 15236
rect 800 14956 59200 14964
rect 800 14556 59120 14956
rect 800 14548 59200 14556
rect 880 14148 59200 14548
rect 800 14140 59200 14148
rect 800 13740 59120 14140
rect 800 13732 59200 13740
rect 880 13332 59200 13732
rect 800 13324 59200 13332
rect 800 12924 59120 13324
rect 800 12916 59200 12924
rect 880 12644 59200 12916
rect 880 12516 59120 12644
rect 800 12244 59120 12516
rect 800 12100 59200 12244
rect 880 11828 59200 12100
rect 880 11700 59120 11828
rect 800 11428 59120 11700
rect 800 11284 59200 11428
rect 880 11148 59200 11284
rect 880 10884 59120 11148
rect 800 10748 59120 10884
rect 800 10468 59200 10748
rect 880 10332 59200 10468
rect 880 10068 59120 10332
rect 800 9932 59120 10068
rect 800 9652 59200 9932
rect 880 9516 59200 9652
rect 880 9252 59120 9516
rect 800 9116 59120 9252
rect 800 8836 59200 9116
rect 880 8436 59120 8836
rect 800 8020 59200 8436
rect 880 7620 59120 8020
rect 800 7340 59200 7620
rect 800 7204 59120 7340
rect 880 6940 59120 7204
rect 880 6804 59200 6940
rect 800 6524 59200 6804
rect 800 6388 59120 6524
rect 880 6124 59120 6388
rect 880 5988 59200 6124
rect 800 5844 59200 5988
rect 800 5572 59120 5844
rect 880 5444 59120 5572
rect 880 5172 59200 5444
rect 800 5028 59200 5172
rect 800 4756 59120 5028
rect 880 4628 59120 4756
rect 880 4356 59200 4628
rect 800 4212 59200 4356
rect 800 3940 59120 4212
rect 880 3812 59120 3940
rect 880 3540 59200 3812
rect 800 3532 59200 3540
rect 800 3132 59120 3532
rect 800 3124 59200 3132
rect 880 2724 59200 3124
rect 800 2716 59200 2724
rect 800 2316 59120 2716
rect 800 2308 59200 2316
rect 880 2036 59200 2308
rect 880 1908 59120 2036
rect 800 1636 59120 1908
rect 800 1492 59200 1636
rect 880 1220 59200 1492
rect 880 1092 59120 1220
rect 800 820 59120 1092
rect 800 676 59200 820
rect 880 540 59200 676
rect 880 511 59120 540
<< metal4 >>
rect 4208 496 4528 57712
rect 19568 496 19888 57712
rect 34928 496 35248 57712
rect 50288 496 50608 57712
<< obsm4 >>
rect 13675 1531 19488 50285
rect 19968 1531 34848 50285
rect 35328 1531 44101 50285
<< labels >>
rlabel metal2 s 542 59200 654 60000 6 active
port 1 nsew signal input
rlabel metal2 s 2934 59200 3046 60000 6 io_in[0]
port 2 nsew signal input
rlabel metal2 s 15170 59200 15282 60000 6 io_in[10]
port 3 nsew signal input
rlabel metal2 s 16366 59200 16478 60000 6 io_in[11]
port 4 nsew signal input
rlabel metal2 s 17654 59200 17766 60000 6 io_in[12]
port 5 nsew signal input
rlabel metal2 s 18850 59200 18962 60000 6 io_in[13]
port 6 nsew signal input
rlabel metal2 s 20046 59200 20158 60000 6 io_in[14]
port 7 nsew signal input
rlabel metal2 s 21334 59200 21446 60000 6 io_in[15]
port 8 nsew signal input
rlabel metal2 s 22530 59200 22642 60000 6 io_in[16]
port 9 nsew signal input
rlabel metal2 s 23726 59200 23838 60000 6 io_in[17]
port 10 nsew signal input
rlabel metal2 s 25014 59200 25126 60000 6 io_in[18]
port 11 nsew signal input
rlabel metal2 s 26210 59200 26322 60000 6 io_in[19]
port 12 nsew signal input
rlabel metal2 s 4130 59200 4242 60000 6 io_in[1]
port 13 nsew signal input
rlabel metal2 s 27406 59200 27518 60000 6 io_in[20]
port 14 nsew signal input
rlabel metal2 s 28694 59200 28806 60000 6 io_in[21]
port 15 nsew signal input
rlabel metal2 s 29890 59200 30002 60000 6 io_in[22]
port 16 nsew signal input
rlabel metal2 s 31086 59200 31198 60000 6 io_in[23]
port 17 nsew signal input
rlabel metal2 s 32282 59200 32394 60000 6 io_in[24]
port 18 nsew signal input
rlabel metal2 s 33570 59200 33682 60000 6 io_in[25]
port 19 nsew signal input
rlabel metal2 s 34766 59200 34878 60000 6 io_in[26]
port 20 nsew signal input
rlabel metal2 s 35962 59200 36074 60000 6 io_in[27]
port 21 nsew signal input
rlabel metal2 s 37250 59200 37362 60000 6 io_in[28]
port 22 nsew signal input
rlabel metal2 s 38446 59200 38558 60000 6 io_in[29]
port 23 nsew signal input
rlabel metal2 s 5418 59200 5530 60000 6 io_in[2]
port 24 nsew signal input
rlabel metal2 s 39642 59200 39754 60000 6 io_in[30]
port 25 nsew signal input
rlabel metal2 s 40930 59200 41042 60000 6 io_in[31]
port 26 nsew signal input
rlabel metal2 s 42126 59200 42238 60000 6 io_in[32]
port 27 nsew signal input
rlabel metal2 s 43322 59200 43434 60000 6 io_in[33]
port 28 nsew signal input
rlabel metal2 s 44610 59200 44722 60000 6 io_in[34]
port 29 nsew signal input
rlabel metal2 s 45806 59200 45918 60000 6 io_in[35]
port 30 nsew signal input
rlabel metal2 s 47002 59200 47114 60000 6 io_in[36]
port 31 nsew signal input
rlabel metal2 s 48198 59200 48310 60000 6 io_in[37]
port 32 nsew signal input
rlabel metal2 s 6614 59200 6726 60000 6 io_in[3]
port 33 nsew signal input
rlabel metal2 s 7810 59200 7922 60000 6 io_in[4]
port 34 nsew signal input
rlabel metal2 s 9098 59200 9210 60000 6 io_in[5]
port 35 nsew signal input
rlabel metal2 s 10294 59200 10406 60000 6 io_in[6]
port 36 nsew signal input
rlabel metal2 s 11490 59200 11602 60000 6 io_in[7]
port 37 nsew signal input
rlabel metal2 s 12778 59200 12890 60000 6 io_in[8]
port 38 nsew signal input
rlabel metal2 s 13974 59200 14086 60000 6 io_in[9]
port 39 nsew signal input
rlabel metal3 s 59200 24428 60000 24668 6 io_oeb[0]
port 40 nsew signal output
rlabel metal3 s 59200 32044 60000 32284 6 io_oeb[10]
port 41 nsew signal output
rlabel metal3 s 59200 32860 60000 33100 6 io_oeb[11]
port 42 nsew signal output
rlabel metal3 s 59200 33540 60000 33780 6 io_oeb[12]
port 43 nsew signal output
rlabel metal3 s 59200 34356 60000 34596 6 io_oeb[13]
port 44 nsew signal output
rlabel metal3 s 59200 35036 60000 35276 6 io_oeb[14]
port 45 nsew signal output
rlabel metal3 s 59200 35852 60000 36092 6 io_oeb[15]
port 46 nsew signal output
rlabel metal3 s 59200 36532 60000 36772 6 io_oeb[16]
port 47 nsew signal output
rlabel metal3 s 59200 37348 60000 37588 6 io_oeb[17]
port 48 nsew signal output
rlabel metal3 s 59200 38164 60000 38404 6 io_oeb[18]
port 49 nsew signal output
rlabel metal3 s 59200 38844 60000 39084 6 io_oeb[19]
port 50 nsew signal output
rlabel metal3 s 59200 25244 60000 25484 6 io_oeb[1]
port 51 nsew signal output
rlabel metal3 s 59200 39660 60000 39900 6 io_oeb[20]
port 52 nsew signal output
rlabel metal3 s 59200 40340 60000 40580 6 io_oeb[21]
port 53 nsew signal output
rlabel metal3 s 59200 41156 60000 41396 6 io_oeb[22]
port 54 nsew signal output
rlabel metal3 s 59200 41972 60000 42212 6 io_oeb[23]
port 55 nsew signal output
rlabel metal3 s 59200 42652 60000 42892 6 io_oeb[24]
port 56 nsew signal output
rlabel metal3 s 59200 43468 60000 43708 6 io_oeb[25]
port 57 nsew signal output
rlabel metal3 s 59200 44148 60000 44388 6 io_oeb[26]
port 58 nsew signal output
rlabel metal3 s 59200 44964 60000 45204 6 io_oeb[27]
port 59 nsew signal output
rlabel metal3 s 59200 45644 60000 45884 6 io_oeb[28]
port 60 nsew signal output
rlabel metal3 s 59200 46460 60000 46700 6 io_oeb[29]
port 61 nsew signal output
rlabel metal3 s 59200 25924 60000 26164 6 io_oeb[2]
port 62 nsew signal output
rlabel metal3 s 59200 47276 60000 47516 6 io_oeb[30]
port 63 nsew signal output
rlabel metal3 s 59200 47956 60000 48196 6 io_oeb[31]
port 64 nsew signal output
rlabel metal3 s 59200 48772 60000 49012 6 io_oeb[32]
port 65 nsew signal output
rlabel metal3 s 59200 49452 60000 49692 6 io_oeb[33]
port 66 nsew signal output
rlabel metal3 s 59200 50268 60000 50508 6 io_oeb[34]
port 67 nsew signal output
rlabel metal3 s 59200 51084 60000 51324 6 io_oeb[35]
port 68 nsew signal output
rlabel metal3 s 59200 51764 60000 52004 6 io_oeb[36]
port 69 nsew signal output
rlabel metal3 s 59200 52580 60000 52820 6 io_oeb[37]
port 70 nsew signal output
rlabel metal3 s 59200 26740 60000 26980 6 io_oeb[3]
port 71 nsew signal output
rlabel metal3 s 59200 27420 60000 27660 6 io_oeb[4]
port 72 nsew signal output
rlabel metal3 s 59200 28236 60000 28476 6 io_oeb[5]
port 73 nsew signal output
rlabel metal3 s 59200 29052 60000 29292 6 io_oeb[6]
port 74 nsew signal output
rlabel metal3 s 59200 29732 60000 29972 6 io_oeb[7]
port 75 nsew signal output
rlabel metal3 s 59200 30548 60000 30788 6 io_oeb[8]
port 76 nsew signal output
rlabel metal3 s 59200 31228 60000 31468 6 io_oeb[9]
port 77 nsew signal output
rlabel metal2 s 49486 59200 49598 60000 6 io_out[0]
port 78 nsew signal output
rlabel metal3 s 59200 54076 60000 54316 6 io_out[10]
port 79 nsew signal output
rlabel metal3 s 59200 54756 60000 54996 6 io_out[11]
port 80 nsew signal output
rlabel metal3 s 59200 55572 60000 55812 6 io_out[12]
port 81 nsew signal output
rlabel metal2 s 8086 0 8198 800 6 io_out[13]
port 82 nsew signal output
rlabel metal3 s 59200 56388 60000 56628 6 io_out[14]
port 83 nsew signal output
rlabel metal2 s 54362 59200 54474 60000 6 io_out[15]
port 84 nsew signal output
rlabel metal2 s 13514 0 13626 800 6 io_out[16]
port 85 nsew signal output
rlabel metal2 s 55558 59200 55670 60000 6 io_out[17]
port 86 nsew signal output
rlabel metal3 s 59200 57068 60000 57308 6 io_out[18]
port 87 nsew signal output
rlabel metal2 s 18942 0 19054 800 6 io_out[19]
port 88 nsew signal output
rlabel metal3 s 59200 53260 60000 53500 6 io_out[1]
port 89 nsew signal output
rlabel metal2 s 24462 0 24574 800 6 io_out[20]
port 90 nsew signal output
rlabel metal2 s 56846 59200 56958 60000 6 io_out[21]
port 91 nsew signal output
rlabel metal2 s 29890 0 30002 800 6 io_out[22]
port 92 nsew signal output
rlabel metal3 s 0 56116 800 56356 6 io_out[23]
port 93 nsew signal output
rlabel metal2 s 35318 0 35430 800 6 io_out[24]
port 94 nsew signal output
rlabel metal2 s 40746 0 40858 800 6 io_out[25]
port 95 nsew signal output
rlabel metal2 s 46266 0 46378 800 6 io_out[26]
port 96 nsew signal output
rlabel metal2 s 58042 59200 58154 60000 6 io_out[27]
port 97 nsew signal output
rlabel metal3 s 59200 57884 60000 58124 6 io_out[28]
port 98 nsew signal output
rlabel metal3 s 0 56932 800 57172 6 io_out[29]
port 99 nsew signal output
rlabel metal2 s 50682 59200 50794 60000 6 io_out[2]
port 100 nsew signal output
rlabel metal3 s 0 57748 800 57988 6 io_out[30]
port 101 nsew signal output
rlabel metal3 s 0 58564 800 58804 6 io_out[31]
port 102 nsew signal output
rlabel metal3 s 0 59380 800 59620 6 io_out[32]
port 103 nsew signal output
rlabel metal3 s 59200 58564 60000 58804 6 io_out[33]
port 104 nsew signal output
rlabel metal2 s 51694 0 51806 800 6 io_out[34]
port 105 nsew signal output
rlabel metal2 s 59238 59200 59350 60000 6 io_out[35]
port 106 nsew signal output
rlabel metal2 s 57122 0 57234 800 6 io_out[36]
port 107 nsew signal output
rlabel metal3 s 59200 59380 60000 59620 6 io_out[37]
port 108 nsew signal output
rlabel metal3 s 0 52852 800 53092 6 io_out[3]
port 109 nsew signal output
rlabel metal3 s 0 53668 800 53908 6 io_out[4]
port 110 nsew signal output
rlabel metal3 s 0 54484 800 54724 6 io_out[5]
port 111 nsew signal output
rlabel metal2 s 51878 59200 51990 60000 6 io_out[6]
port 112 nsew signal output
rlabel metal2 s 53166 59200 53278 60000 6 io_out[7]
port 113 nsew signal output
rlabel metal3 s 0 55300 800 55540 6 io_out[8]
port 114 nsew signal output
rlabel metal2 s 2658 0 2770 800 6 io_out[9]
port 115 nsew signal output
rlabel metal3 s 0 356 800 596 6 la1_data_in[0]
port 116 nsew signal input
rlabel metal3 s 0 8516 800 8756 6 la1_data_in[10]
port 117 nsew signal input
rlabel metal3 s 0 9332 800 9572 6 la1_data_in[11]
port 118 nsew signal input
rlabel metal3 s 0 10148 800 10388 6 la1_data_in[12]
port 119 nsew signal input
rlabel metal3 s 0 10964 800 11204 6 la1_data_in[13]
port 120 nsew signal input
rlabel metal3 s 0 11780 800 12020 6 la1_data_in[14]
port 121 nsew signal input
rlabel metal3 s 0 12596 800 12836 6 la1_data_in[15]
port 122 nsew signal input
rlabel metal3 s 0 13412 800 13652 6 la1_data_in[16]
port 123 nsew signal input
rlabel metal3 s 0 14228 800 14468 6 la1_data_in[17]
port 124 nsew signal input
rlabel metal3 s 0 15044 800 15284 6 la1_data_in[18]
port 125 nsew signal input
rlabel metal3 s 0 15860 800 16100 6 la1_data_in[19]
port 126 nsew signal input
rlabel metal3 s 0 1172 800 1412 6 la1_data_in[1]
port 127 nsew signal input
rlabel metal3 s 0 16676 800 16916 6 la1_data_in[20]
port 128 nsew signal input
rlabel metal3 s 0 17492 800 17732 6 la1_data_in[21]
port 129 nsew signal input
rlabel metal3 s 0 18308 800 18548 6 la1_data_in[22]
port 130 nsew signal input
rlabel metal3 s 0 19124 800 19364 6 la1_data_in[23]
port 131 nsew signal input
rlabel metal3 s 0 19940 800 20180 6 la1_data_in[24]
port 132 nsew signal input
rlabel metal3 s 0 20892 800 21132 6 la1_data_in[25]
port 133 nsew signal input
rlabel metal3 s 0 21708 800 21948 6 la1_data_in[26]
port 134 nsew signal input
rlabel metal3 s 0 22524 800 22764 6 la1_data_in[27]
port 135 nsew signal input
rlabel metal3 s 0 23340 800 23580 6 la1_data_in[28]
port 136 nsew signal input
rlabel metal3 s 0 24156 800 24396 6 la1_data_in[29]
port 137 nsew signal input
rlabel metal3 s 0 1988 800 2228 6 la1_data_in[2]
port 138 nsew signal input
rlabel metal3 s 0 24972 800 25212 6 la1_data_in[30]
port 139 nsew signal input
rlabel metal3 s 0 25788 800 26028 6 la1_data_in[31]
port 140 nsew signal input
rlabel metal3 s 0 2804 800 3044 6 la1_data_in[3]
port 141 nsew signal input
rlabel metal3 s 0 3620 800 3860 6 la1_data_in[4]
port 142 nsew signal input
rlabel metal3 s 0 4436 800 4676 6 la1_data_in[5]
port 143 nsew signal input
rlabel metal3 s 0 5252 800 5492 6 la1_data_in[6]
port 144 nsew signal input
rlabel metal3 s 0 6068 800 6308 6 la1_data_in[7]
port 145 nsew signal input
rlabel metal3 s 0 6884 800 7124 6 la1_data_in[8]
port 146 nsew signal input
rlabel metal3 s 0 7700 800 7940 6 la1_data_in[9]
port 147 nsew signal input
rlabel metal3 s 0 26604 800 26844 6 la1_data_out[0]
port 148 nsew signal output
rlabel metal3 s 0 34764 800 35004 6 la1_data_out[10]
port 149 nsew signal output
rlabel metal3 s 0 35580 800 35820 6 la1_data_out[11]
port 150 nsew signal output
rlabel metal3 s 0 36396 800 36636 6 la1_data_out[12]
port 151 nsew signal output
rlabel metal3 s 0 37212 800 37452 6 la1_data_out[13]
port 152 nsew signal output
rlabel metal3 s 0 38028 800 38268 6 la1_data_out[14]
port 153 nsew signal output
rlabel metal3 s 0 38844 800 39084 6 la1_data_out[15]
port 154 nsew signal output
rlabel metal3 s 0 39660 800 39900 6 la1_data_out[16]
port 155 nsew signal output
rlabel metal3 s 0 40612 800 40852 6 la1_data_out[17]
port 156 nsew signal output
rlabel metal3 s 0 41428 800 41668 6 la1_data_out[18]
port 157 nsew signal output
rlabel metal3 s 0 42244 800 42484 6 la1_data_out[19]
port 158 nsew signal output
rlabel metal3 s 0 27420 800 27660 6 la1_data_out[1]
port 159 nsew signal output
rlabel metal3 s 0 43060 800 43300 6 la1_data_out[20]
port 160 nsew signal output
rlabel metal3 s 0 43876 800 44116 6 la1_data_out[21]
port 161 nsew signal output
rlabel metal3 s 0 44692 800 44932 6 la1_data_out[22]
port 162 nsew signal output
rlabel metal3 s 0 45508 800 45748 6 la1_data_out[23]
port 163 nsew signal output
rlabel metal3 s 0 46324 800 46564 6 la1_data_out[24]
port 164 nsew signal output
rlabel metal3 s 0 47140 800 47380 6 la1_data_out[25]
port 165 nsew signal output
rlabel metal3 s 0 47956 800 48196 6 la1_data_out[26]
port 166 nsew signal output
rlabel metal3 s 0 48772 800 49012 6 la1_data_out[27]
port 167 nsew signal output
rlabel metal3 s 0 49588 800 49828 6 la1_data_out[28]
port 168 nsew signal output
rlabel metal3 s 0 50404 800 50644 6 la1_data_out[29]
port 169 nsew signal output
rlabel metal3 s 0 28236 800 28476 6 la1_data_out[2]
port 170 nsew signal output
rlabel metal3 s 0 51220 800 51460 6 la1_data_out[30]
port 171 nsew signal output
rlabel metal3 s 0 52036 800 52276 6 la1_data_out[31]
port 172 nsew signal output
rlabel metal3 s 0 29052 800 29292 6 la1_data_out[3]
port 173 nsew signal output
rlabel metal3 s 0 29868 800 30108 6 la1_data_out[4]
port 174 nsew signal output
rlabel metal3 s 0 30684 800 30924 6 la1_data_out[5]
port 175 nsew signal output
rlabel metal3 s 0 31500 800 31740 6 la1_data_out[6]
port 176 nsew signal output
rlabel metal3 s 0 32316 800 32556 6 la1_data_out[7]
port 177 nsew signal output
rlabel metal3 s 0 33132 800 33372 6 la1_data_out[8]
port 178 nsew signal output
rlabel metal3 s 0 33948 800 34188 6 la1_data_out[9]
port 179 nsew signal output
rlabel metal3 s 59200 220 60000 460 6 la1_oenb[0]
port 180 nsew signal input
rlabel metal3 s 59200 7700 60000 7940 6 la1_oenb[10]
port 181 nsew signal input
rlabel metal3 s 59200 8516 60000 8756 6 la1_oenb[11]
port 182 nsew signal input
rlabel metal3 s 59200 9196 60000 9436 6 la1_oenb[12]
port 183 nsew signal input
rlabel metal3 s 59200 10012 60000 10252 6 la1_oenb[13]
port 184 nsew signal input
rlabel metal3 s 59200 10828 60000 11068 6 la1_oenb[14]
port 185 nsew signal input
rlabel metal3 s 59200 11508 60000 11748 6 la1_oenb[15]
port 186 nsew signal input
rlabel metal3 s 59200 12324 60000 12564 6 la1_oenb[16]
port 187 nsew signal input
rlabel metal3 s 59200 13004 60000 13244 6 la1_oenb[17]
port 188 nsew signal input
rlabel metal3 s 59200 13820 60000 14060 6 la1_oenb[18]
port 189 nsew signal input
rlabel metal3 s 59200 14636 60000 14876 6 la1_oenb[19]
port 190 nsew signal input
rlabel metal3 s 59200 900 60000 1140 6 la1_oenb[1]
port 191 nsew signal input
rlabel metal3 s 59200 15316 60000 15556 6 la1_oenb[20]
port 192 nsew signal input
rlabel metal3 s 59200 16132 60000 16372 6 la1_oenb[21]
port 193 nsew signal input
rlabel metal3 s 59200 16812 60000 17052 6 la1_oenb[22]
port 194 nsew signal input
rlabel metal3 s 59200 17628 60000 17868 6 la1_oenb[23]
port 195 nsew signal input
rlabel metal3 s 59200 18308 60000 18548 6 la1_oenb[24]
port 196 nsew signal input
rlabel metal3 s 59200 19124 60000 19364 6 la1_oenb[25]
port 197 nsew signal input
rlabel metal3 s 59200 19940 60000 20180 6 la1_oenb[26]
port 198 nsew signal input
rlabel metal3 s 59200 20620 60000 20860 6 la1_oenb[27]
port 199 nsew signal input
rlabel metal3 s 59200 21436 60000 21676 6 la1_oenb[28]
port 200 nsew signal input
rlabel metal3 s 59200 22116 60000 22356 6 la1_oenb[29]
port 201 nsew signal input
rlabel metal3 s 59200 1716 60000 1956 6 la1_oenb[2]
port 202 nsew signal input
rlabel metal3 s 59200 22932 60000 23172 6 la1_oenb[30]
port 203 nsew signal input
rlabel metal3 s 59200 23748 60000 23988 6 la1_oenb[31]
port 204 nsew signal input
rlabel metal3 s 59200 2396 60000 2636 6 la1_oenb[3]
port 205 nsew signal input
rlabel metal3 s 59200 3212 60000 3452 6 la1_oenb[4]
port 206 nsew signal input
rlabel metal3 s 59200 3892 60000 4132 6 la1_oenb[5]
port 207 nsew signal input
rlabel metal3 s 59200 4708 60000 4948 6 la1_oenb[6]
port 208 nsew signal input
rlabel metal3 s 59200 5524 60000 5764 6 la1_oenb[7]
port 209 nsew signal input
rlabel metal3 s 59200 6204 60000 6444 6 la1_oenb[8]
port 210 nsew signal input
rlabel metal3 s 59200 7020 60000 7260 6 la1_oenb[9]
port 211 nsew signal input
rlabel metal4 s 4208 496 4528 57712 6 vccd1
port 212 nsew power input
rlabel metal4 s 34928 496 35248 57712 6 vccd1
port 212 nsew power input
rlabel metal4 s 19568 496 19888 57712 6 vssd1
port 213 nsew ground input
rlabel metal4 s 50288 496 50608 57712 6 vssd1
port 213 nsew ground input
rlabel metal2 s 1738 59200 1850 60000 6 wb_clk_i
port 214 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 60000 60000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 12605898
string GDS_FILE /openlane/designs/wrapped-vgademo-on-fpga/runs/RUN_2022.03.20_08.41.27/results/finishing/wrapped_vgademo_on_fpga.magic.gds
string GDS_START 1090208
<< end >>

