magic
tech sky130A
magscale 1 2
timestamp 1647739228
<< obsli1 >>
rect 1104 527 58880 53329
<< obsm1 >>
rect 382 496 59602 54392
<< metal2 >>
rect 358 55200 470 56000
rect 1094 55200 1206 56000
rect 1830 55200 1942 56000
rect 2658 55200 2770 56000
rect 3394 55200 3506 56000
rect 4130 55200 4242 56000
rect 4958 55200 5070 56000
rect 5694 55200 5806 56000
rect 6430 55200 6542 56000
rect 7258 55200 7370 56000
rect 7994 55200 8106 56000
rect 8730 55200 8842 56000
rect 9558 55200 9670 56000
rect 10294 55200 10406 56000
rect 11122 55200 11234 56000
rect 11858 55200 11970 56000
rect 12594 55200 12706 56000
rect 13422 55200 13534 56000
rect 14158 55200 14270 56000
rect 14894 55200 15006 56000
rect 15722 55200 15834 56000
rect 16458 55200 16570 56000
rect 17194 55200 17306 56000
rect 18022 55200 18134 56000
rect 18758 55200 18870 56000
rect 19494 55200 19606 56000
rect 20322 55200 20434 56000
rect 21058 55200 21170 56000
rect 21886 55200 21998 56000
rect 22622 55200 22734 56000
rect 23358 55200 23470 56000
rect 24186 55200 24298 56000
rect 24922 55200 25034 56000
rect 25658 55200 25770 56000
rect 26486 55200 26598 56000
rect 27222 55200 27334 56000
rect 27958 55200 28070 56000
rect 28786 55200 28898 56000
rect 29522 55200 29634 56000
rect 30350 55200 30462 56000
rect 31086 55200 31198 56000
rect 31822 55200 31934 56000
rect 32650 55200 32762 56000
rect 33386 55200 33498 56000
rect 34122 55200 34234 56000
rect 34950 55200 35062 56000
rect 35686 55200 35798 56000
rect 36422 55200 36534 56000
rect 37250 55200 37362 56000
rect 37986 55200 38098 56000
rect 38722 55200 38834 56000
rect 39550 55200 39662 56000
rect 40286 55200 40398 56000
rect 41114 55200 41226 56000
rect 41850 55200 41962 56000
rect 42586 55200 42698 56000
rect 43414 55200 43526 56000
rect 44150 55200 44262 56000
rect 44886 55200 44998 56000
rect 45714 55200 45826 56000
rect 46450 55200 46562 56000
rect 47186 55200 47298 56000
rect 48014 55200 48126 56000
rect 48750 55200 48862 56000
rect 49486 55200 49598 56000
rect 50314 55200 50426 56000
rect 51050 55200 51162 56000
rect 51878 55200 51990 56000
rect 52614 55200 52726 56000
rect 53350 55200 53462 56000
rect 54178 55200 54290 56000
rect 54914 55200 55026 56000
rect 55650 55200 55762 56000
rect 56478 55200 56590 56000
rect 57214 55200 57326 56000
rect 57950 55200 58062 56000
rect 58778 55200 58890 56000
rect 59514 55200 59626 56000
<< obsm2 >>
rect 526 55144 1038 55593
rect 1262 55144 1774 55593
rect 1998 55144 2602 55593
rect 2826 55144 3338 55593
rect 3562 55144 4074 55593
rect 4298 55144 4902 55593
rect 5126 55144 5638 55593
rect 5862 55144 6374 55593
rect 6598 55144 7202 55593
rect 7426 55144 7938 55593
rect 8162 55144 8674 55593
rect 8898 55144 9502 55593
rect 9726 55144 10238 55593
rect 10462 55144 11066 55593
rect 11290 55144 11802 55593
rect 12026 55144 12538 55593
rect 12762 55144 13366 55593
rect 13590 55144 14102 55593
rect 14326 55144 14838 55593
rect 15062 55144 15666 55593
rect 15890 55144 16402 55593
rect 16626 55144 17138 55593
rect 17362 55144 17966 55593
rect 18190 55144 18702 55593
rect 18926 55144 19438 55593
rect 19662 55144 20266 55593
rect 20490 55144 21002 55593
rect 21226 55144 21830 55593
rect 22054 55144 22566 55593
rect 22790 55144 23302 55593
rect 23526 55144 24130 55593
rect 24354 55144 24866 55593
rect 25090 55144 25602 55593
rect 25826 55144 26430 55593
rect 26654 55144 27166 55593
rect 27390 55144 27902 55593
rect 28126 55144 28730 55593
rect 28954 55144 29466 55593
rect 29690 55144 30294 55593
rect 30518 55144 31030 55593
rect 31254 55144 31766 55593
rect 31990 55144 32594 55593
rect 32818 55144 33330 55593
rect 33554 55144 34066 55593
rect 34290 55144 34894 55593
rect 35118 55144 35630 55593
rect 35854 55144 36366 55593
rect 36590 55144 37194 55593
rect 37418 55144 37930 55593
rect 38154 55144 38666 55593
rect 38890 55144 39494 55593
rect 39718 55144 40230 55593
rect 40454 55144 41058 55593
rect 41282 55144 41794 55593
rect 42018 55144 42530 55593
rect 42754 55144 43358 55593
rect 43582 55144 44094 55593
rect 44318 55144 44830 55593
rect 45054 55144 45658 55593
rect 45882 55144 46394 55593
rect 46618 55144 47130 55593
rect 47354 55144 47958 55593
rect 48182 55144 48694 55593
rect 48918 55144 49430 55593
rect 49654 55144 50258 55593
rect 50482 55144 50994 55593
rect 51218 55144 51822 55593
rect 52046 55144 52558 55593
rect 52782 55144 53294 55593
rect 53518 55144 54122 55593
rect 54346 55144 54858 55593
rect 55082 55144 55594 55593
rect 55818 55144 56422 55593
rect 56646 55144 57158 55593
rect 57382 55144 57894 55593
rect 58118 55144 58722 55593
rect 58946 55144 59458 55593
rect 388 496 59596 55144
<< metal3 >>
rect 0 55436 800 55676
rect 59200 55436 60000 55676
rect 0 54620 800 54860
rect 59200 54620 60000 54860
rect 0 53668 800 53908
rect 59200 53804 60000 54044
rect 0 52852 800 53092
rect 59200 52988 60000 53228
rect 0 51900 800 52140
rect 59200 52172 60000 52412
rect 0 51084 800 51324
rect 59200 51356 60000 51596
rect 59200 50540 60000 50780
rect 0 50132 800 50372
rect 59200 49724 60000 49964
rect 0 49316 800 49556
rect 59200 49044 60000 49284
rect 0 48500 800 48740
rect 59200 48228 60000 48468
rect 0 47548 800 47788
rect 59200 47412 60000 47652
rect 0 46732 800 46972
rect 59200 46596 60000 46836
rect 0 45780 800 46020
rect 59200 45780 60000 46020
rect 0 44964 800 45204
rect 59200 44964 60000 45204
rect 0 44012 800 44252
rect 59200 44148 60000 44388
rect 0 43196 800 43436
rect 59200 43332 60000 43572
rect 0 42380 800 42620
rect 59200 42516 60000 42756
rect 59200 41836 60000 42076
rect 0 41428 800 41668
rect 59200 41020 60000 41260
rect 0 40612 800 40852
rect 59200 40204 60000 40444
rect 0 39660 800 39900
rect 59200 39388 60000 39628
rect 0 38844 800 39084
rect 59200 38572 60000 38812
rect 0 37892 800 38132
rect 59200 37756 60000 37996
rect 0 37076 800 37316
rect 59200 36940 60000 37180
rect 0 36124 800 36364
rect 59200 36124 60000 36364
rect 0 35308 800 35548
rect 59200 35308 60000 35548
rect 0 34492 800 34732
rect 59200 34628 60000 34868
rect 0 33540 800 33780
rect 59200 33812 60000 34052
rect 0 32724 800 32964
rect 59200 32996 60000 33236
rect 59200 32180 60000 32420
rect 0 31772 800 32012
rect 59200 31364 60000 31604
rect 0 30956 800 31196
rect 59200 30548 60000 30788
rect 0 30004 800 30244
rect 59200 29732 60000 29972
rect 0 29188 800 29428
rect 59200 28916 60000 29156
rect 0 28372 800 28612
rect 59200 28236 60000 28476
rect 0 27420 800 27660
rect 59200 27420 60000 27660
rect 0 26604 800 26844
rect 59200 26604 60000 26844
rect 0 25652 800 25892
rect 59200 25788 60000 26028
rect 0 24836 800 25076
rect 59200 24972 60000 25212
rect 0 23884 800 24124
rect 59200 24156 60000 24396
rect 0 23068 800 23308
rect 59200 23340 60000 23580
rect 59200 22524 60000 22764
rect 0 22116 800 22356
rect 59200 21708 60000 21948
rect 0 21300 800 21540
rect 59200 21028 60000 21268
rect 0 20484 800 20724
rect 59200 20212 60000 20452
rect 0 19532 800 19772
rect 59200 19396 60000 19636
rect 0 18716 800 18956
rect 59200 18580 60000 18820
rect 0 17764 800 18004
rect 59200 17764 60000 18004
rect 0 16948 800 17188
rect 59200 16948 60000 17188
rect 0 15996 800 16236
rect 59200 16132 60000 16372
rect 0 15180 800 15420
rect 59200 15316 60000 15556
rect 0 14364 800 14604
rect 59200 14500 60000 14740
rect 59200 13820 60000 14060
rect 0 13412 800 13652
rect 59200 13004 60000 13244
rect 0 12596 800 12836
rect 59200 12188 60000 12428
rect 0 11644 800 11884
rect 59200 11372 60000 11612
rect 0 10828 800 11068
rect 59200 10556 60000 10796
rect 0 9876 800 10116
rect 59200 9740 60000 9980
rect 0 9060 800 9300
rect 59200 8924 60000 9164
rect 0 8108 800 8348
rect 59200 8108 60000 8348
rect 0 7292 800 7532
rect 59200 7292 60000 7532
rect 0 6476 800 6716
rect 59200 6612 60000 6852
rect 0 5524 800 5764
rect 59200 5796 60000 6036
rect 0 4708 800 4948
rect 59200 4980 60000 5220
rect 59200 4164 60000 4404
rect 0 3756 800 3996
rect 59200 3348 60000 3588
rect 0 2940 800 3180
rect 59200 2532 60000 2772
rect 0 1988 800 2228
rect 59200 1716 60000 1956
rect 0 1172 800 1412
rect 59200 900 60000 1140
rect 0 356 800 596
rect 59200 220 60000 460
<< obsm3 >>
rect 880 55356 59120 55589
rect 800 54940 59200 55356
rect 880 54540 59120 54940
rect 800 54124 59200 54540
rect 800 53988 59120 54124
rect 880 53724 59120 53988
rect 880 53588 59200 53724
rect 800 53308 59200 53588
rect 800 53172 59120 53308
rect 880 52908 59120 53172
rect 880 52772 59200 52908
rect 800 52492 59200 52772
rect 800 52220 59120 52492
rect 880 52092 59120 52220
rect 880 51820 59200 52092
rect 800 51676 59200 51820
rect 800 51404 59120 51676
rect 880 51276 59120 51404
rect 880 51004 59200 51276
rect 800 50860 59200 51004
rect 800 50460 59120 50860
rect 800 50452 59200 50460
rect 880 50052 59200 50452
rect 800 50044 59200 50052
rect 800 49644 59120 50044
rect 800 49636 59200 49644
rect 880 49364 59200 49636
rect 880 49236 59120 49364
rect 800 48964 59120 49236
rect 800 48820 59200 48964
rect 880 48548 59200 48820
rect 880 48420 59120 48548
rect 800 48148 59120 48420
rect 800 47868 59200 48148
rect 880 47732 59200 47868
rect 880 47468 59120 47732
rect 800 47332 59120 47468
rect 800 47052 59200 47332
rect 880 46916 59200 47052
rect 880 46652 59120 46916
rect 800 46516 59120 46652
rect 800 46100 59200 46516
rect 880 45700 59120 46100
rect 800 45284 59200 45700
rect 880 44884 59120 45284
rect 800 44468 59200 44884
rect 800 44332 59120 44468
rect 880 44068 59120 44332
rect 880 43932 59200 44068
rect 800 43652 59200 43932
rect 800 43516 59120 43652
rect 880 43252 59120 43516
rect 880 43116 59200 43252
rect 800 42836 59200 43116
rect 800 42700 59120 42836
rect 880 42436 59120 42700
rect 880 42300 59200 42436
rect 800 42156 59200 42300
rect 800 41756 59120 42156
rect 800 41748 59200 41756
rect 880 41348 59200 41748
rect 800 41340 59200 41348
rect 800 40940 59120 41340
rect 800 40932 59200 40940
rect 880 40532 59200 40932
rect 800 40524 59200 40532
rect 800 40124 59120 40524
rect 800 39980 59200 40124
rect 880 39708 59200 39980
rect 880 39580 59120 39708
rect 800 39308 59120 39580
rect 800 39164 59200 39308
rect 880 38892 59200 39164
rect 880 38764 59120 38892
rect 800 38492 59120 38764
rect 800 38212 59200 38492
rect 880 38076 59200 38212
rect 880 37812 59120 38076
rect 800 37676 59120 37812
rect 800 37396 59200 37676
rect 880 37260 59200 37396
rect 880 36996 59120 37260
rect 800 36860 59120 36996
rect 800 36444 59200 36860
rect 880 36044 59120 36444
rect 800 35628 59200 36044
rect 880 35228 59120 35628
rect 800 34948 59200 35228
rect 800 34812 59120 34948
rect 880 34548 59120 34812
rect 880 34412 59200 34548
rect 800 34132 59200 34412
rect 800 33860 59120 34132
rect 880 33732 59120 33860
rect 880 33460 59200 33732
rect 800 33316 59200 33460
rect 800 33044 59120 33316
rect 880 32916 59120 33044
rect 880 32644 59200 32916
rect 800 32500 59200 32644
rect 800 32100 59120 32500
rect 800 32092 59200 32100
rect 880 31692 59200 32092
rect 800 31684 59200 31692
rect 800 31284 59120 31684
rect 800 31276 59200 31284
rect 880 30876 59200 31276
rect 800 30868 59200 30876
rect 800 30468 59120 30868
rect 800 30324 59200 30468
rect 880 30052 59200 30324
rect 880 29924 59120 30052
rect 800 29652 59120 29924
rect 800 29508 59200 29652
rect 880 29236 59200 29508
rect 880 29108 59120 29236
rect 800 28836 59120 29108
rect 800 28692 59200 28836
rect 880 28556 59200 28692
rect 880 28292 59120 28556
rect 800 28156 59120 28292
rect 800 27740 59200 28156
rect 880 27340 59120 27740
rect 800 26924 59200 27340
rect 880 26524 59120 26924
rect 800 26108 59200 26524
rect 800 25972 59120 26108
rect 880 25708 59120 25972
rect 880 25572 59200 25708
rect 800 25292 59200 25572
rect 800 25156 59120 25292
rect 880 24892 59120 25156
rect 880 24756 59200 24892
rect 800 24476 59200 24756
rect 800 24204 59120 24476
rect 880 24076 59120 24204
rect 880 23804 59200 24076
rect 800 23660 59200 23804
rect 800 23388 59120 23660
rect 880 23260 59120 23388
rect 880 22988 59200 23260
rect 800 22844 59200 22988
rect 800 22444 59120 22844
rect 800 22436 59200 22444
rect 880 22036 59200 22436
rect 800 22028 59200 22036
rect 800 21628 59120 22028
rect 800 21620 59200 21628
rect 880 21348 59200 21620
rect 880 21220 59120 21348
rect 800 20948 59120 21220
rect 800 20804 59200 20948
rect 880 20532 59200 20804
rect 880 20404 59120 20532
rect 800 20132 59120 20404
rect 800 19852 59200 20132
rect 880 19716 59200 19852
rect 880 19452 59120 19716
rect 800 19316 59120 19452
rect 800 19036 59200 19316
rect 880 18900 59200 19036
rect 880 18636 59120 18900
rect 800 18500 59120 18636
rect 800 18084 59200 18500
rect 880 17684 59120 18084
rect 800 17268 59200 17684
rect 880 16868 59120 17268
rect 800 16452 59200 16868
rect 800 16316 59120 16452
rect 880 16052 59120 16316
rect 880 15916 59200 16052
rect 800 15636 59200 15916
rect 800 15500 59120 15636
rect 880 15236 59120 15500
rect 880 15100 59200 15236
rect 800 14820 59200 15100
rect 800 14684 59120 14820
rect 880 14420 59120 14684
rect 880 14284 59200 14420
rect 800 14140 59200 14284
rect 800 13740 59120 14140
rect 800 13732 59200 13740
rect 880 13332 59200 13732
rect 800 13324 59200 13332
rect 800 12924 59120 13324
rect 800 12916 59200 12924
rect 880 12516 59200 12916
rect 800 12508 59200 12516
rect 800 12108 59120 12508
rect 800 11964 59200 12108
rect 880 11692 59200 11964
rect 880 11564 59120 11692
rect 800 11292 59120 11564
rect 800 11148 59200 11292
rect 880 10876 59200 11148
rect 880 10748 59120 10876
rect 800 10476 59120 10748
rect 800 10196 59200 10476
rect 880 10060 59200 10196
rect 880 9796 59120 10060
rect 800 9660 59120 9796
rect 800 9380 59200 9660
rect 880 9244 59200 9380
rect 880 8980 59120 9244
rect 800 8844 59120 8980
rect 800 8428 59200 8844
rect 880 8028 59120 8428
rect 800 7612 59200 8028
rect 880 7212 59120 7612
rect 800 6932 59200 7212
rect 800 6796 59120 6932
rect 880 6532 59120 6796
rect 880 6396 59200 6532
rect 800 6116 59200 6396
rect 800 5844 59120 6116
rect 880 5716 59120 5844
rect 880 5444 59200 5716
rect 800 5300 59200 5444
rect 800 5028 59120 5300
rect 880 4900 59120 5028
rect 880 4628 59200 4900
rect 800 4484 59200 4628
rect 800 4084 59120 4484
rect 800 4076 59200 4084
rect 880 3676 59200 4076
rect 800 3668 59200 3676
rect 800 3268 59120 3668
rect 800 3260 59200 3268
rect 880 2860 59200 3260
rect 800 2852 59200 2860
rect 800 2452 59120 2852
rect 800 2308 59200 2452
rect 880 2036 59200 2308
rect 880 1908 59120 2036
rect 800 1636 59120 1908
rect 800 1492 59200 1636
rect 880 1220 59200 1492
rect 880 1092 59120 1220
rect 800 820 59120 1092
rect 800 676 59200 820
rect 880 540 59200 676
rect 880 511 59120 540
<< metal4 >>
rect 4208 496 4528 53360
rect 19568 496 19888 53360
rect 34928 496 35248 53360
rect 50288 496 50608 53360
<< obsm4 >>
rect 1531 53440 56245 54229
rect 1531 14315 4128 53440
rect 4608 14315 19488 53440
rect 19968 14315 34848 53440
rect 35328 14315 50208 53440
rect 50688 14315 56245 53440
<< labels >>
rlabel metal2 s 358 55200 470 56000 6 active
port 1 nsew signal input
rlabel metal2 s 1830 55200 1942 56000 6 io_in[0]
port 2 nsew signal input
rlabel metal2 s 9558 55200 9670 56000 6 io_in[10]
port 3 nsew signal input
rlabel metal2 s 10294 55200 10406 56000 6 io_in[11]
port 4 nsew signal input
rlabel metal2 s 11122 55200 11234 56000 6 io_in[12]
port 5 nsew signal input
rlabel metal2 s 11858 55200 11970 56000 6 io_in[13]
port 6 nsew signal input
rlabel metal2 s 12594 55200 12706 56000 6 io_in[14]
port 7 nsew signal input
rlabel metal2 s 13422 55200 13534 56000 6 io_in[15]
port 8 nsew signal input
rlabel metal2 s 14158 55200 14270 56000 6 io_in[16]
port 9 nsew signal input
rlabel metal2 s 14894 55200 15006 56000 6 io_in[17]
port 10 nsew signal input
rlabel metal2 s 15722 55200 15834 56000 6 io_in[18]
port 11 nsew signal input
rlabel metal2 s 16458 55200 16570 56000 6 io_in[19]
port 12 nsew signal input
rlabel metal2 s 2658 55200 2770 56000 6 io_in[1]
port 13 nsew signal input
rlabel metal2 s 17194 55200 17306 56000 6 io_in[20]
port 14 nsew signal input
rlabel metal2 s 18022 55200 18134 56000 6 io_in[21]
port 15 nsew signal input
rlabel metal2 s 18758 55200 18870 56000 6 io_in[22]
port 16 nsew signal input
rlabel metal2 s 19494 55200 19606 56000 6 io_in[23]
port 17 nsew signal input
rlabel metal2 s 20322 55200 20434 56000 6 io_in[24]
port 18 nsew signal input
rlabel metal2 s 21058 55200 21170 56000 6 io_in[25]
port 19 nsew signal input
rlabel metal2 s 21886 55200 21998 56000 6 io_in[26]
port 20 nsew signal input
rlabel metal2 s 22622 55200 22734 56000 6 io_in[27]
port 21 nsew signal input
rlabel metal2 s 23358 55200 23470 56000 6 io_in[28]
port 22 nsew signal input
rlabel metal2 s 24186 55200 24298 56000 6 io_in[29]
port 23 nsew signal input
rlabel metal2 s 3394 55200 3506 56000 6 io_in[2]
port 24 nsew signal input
rlabel metal2 s 24922 55200 25034 56000 6 io_in[30]
port 25 nsew signal input
rlabel metal2 s 25658 55200 25770 56000 6 io_in[31]
port 26 nsew signal input
rlabel metal2 s 26486 55200 26598 56000 6 io_in[32]
port 27 nsew signal input
rlabel metal2 s 27222 55200 27334 56000 6 io_in[33]
port 28 nsew signal input
rlabel metal2 s 27958 55200 28070 56000 6 io_in[34]
port 29 nsew signal input
rlabel metal2 s 28786 55200 28898 56000 6 io_in[35]
port 30 nsew signal input
rlabel metal2 s 29522 55200 29634 56000 6 io_in[36]
port 31 nsew signal input
rlabel metal2 s 30350 55200 30462 56000 6 io_in[37]
port 32 nsew signal input
rlabel metal2 s 4130 55200 4242 56000 6 io_in[3]
port 33 nsew signal input
rlabel metal2 s 4958 55200 5070 56000 6 io_in[4]
port 34 nsew signal input
rlabel metal2 s 5694 55200 5806 56000 6 io_in[5]
port 35 nsew signal input
rlabel metal2 s 6430 55200 6542 56000 6 io_in[6]
port 36 nsew signal input
rlabel metal2 s 7258 55200 7370 56000 6 io_in[7]
port 37 nsew signal input
rlabel metal2 s 7994 55200 8106 56000 6 io_in[8]
port 38 nsew signal input
rlabel metal2 s 8730 55200 8842 56000 6 io_in[9]
port 39 nsew signal input
rlabel metal3 s 59200 25788 60000 26028 6 io_oeb[0]
port 40 nsew signal output
rlabel metal3 s 59200 33812 60000 34052 6 io_oeb[10]
port 41 nsew signal output
rlabel metal3 s 59200 34628 60000 34868 6 io_oeb[11]
port 42 nsew signal output
rlabel metal3 s 59200 35308 60000 35548 6 io_oeb[12]
port 43 nsew signal output
rlabel metal3 s 59200 36124 60000 36364 6 io_oeb[13]
port 44 nsew signal output
rlabel metal3 s 59200 36940 60000 37180 6 io_oeb[14]
port 45 nsew signal output
rlabel metal3 s 59200 37756 60000 37996 6 io_oeb[15]
port 46 nsew signal output
rlabel metal3 s 59200 38572 60000 38812 6 io_oeb[16]
port 47 nsew signal output
rlabel metal3 s 59200 39388 60000 39628 6 io_oeb[17]
port 48 nsew signal output
rlabel metal3 s 59200 40204 60000 40444 6 io_oeb[18]
port 49 nsew signal output
rlabel metal3 s 59200 41020 60000 41260 6 io_oeb[19]
port 50 nsew signal output
rlabel metal3 s 59200 26604 60000 26844 6 io_oeb[1]
port 51 nsew signal output
rlabel metal3 s 59200 41836 60000 42076 6 io_oeb[20]
port 52 nsew signal output
rlabel metal3 s 59200 42516 60000 42756 6 io_oeb[21]
port 53 nsew signal output
rlabel metal3 s 59200 43332 60000 43572 6 io_oeb[22]
port 54 nsew signal output
rlabel metal3 s 59200 44148 60000 44388 6 io_oeb[23]
port 55 nsew signal output
rlabel metal3 s 59200 44964 60000 45204 6 io_oeb[24]
port 56 nsew signal output
rlabel metal3 s 59200 45780 60000 46020 6 io_oeb[25]
port 57 nsew signal output
rlabel metal3 s 59200 46596 60000 46836 6 io_oeb[26]
port 58 nsew signal output
rlabel metal3 s 59200 47412 60000 47652 6 io_oeb[27]
port 59 nsew signal output
rlabel metal3 s 59200 48228 60000 48468 6 io_oeb[28]
port 60 nsew signal output
rlabel metal3 s 59200 49044 60000 49284 6 io_oeb[29]
port 61 nsew signal output
rlabel metal3 s 59200 27420 60000 27660 6 io_oeb[2]
port 62 nsew signal output
rlabel metal3 s 59200 49724 60000 49964 6 io_oeb[30]
port 63 nsew signal output
rlabel metal3 s 59200 50540 60000 50780 6 io_oeb[31]
port 64 nsew signal output
rlabel metal3 s 59200 51356 60000 51596 6 io_oeb[32]
port 65 nsew signal output
rlabel metal3 s 59200 52172 60000 52412 6 io_oeb[33]
port 66 nsew signal output
rlabel metal3 s 59200 52988 60000 53228 6 io_oeb[34]
port 67 nsew signal output
rlabel metal3 s 59200 53804 60000 54044 6 io_oeb[35]
port 68 nsew signal output
rlabel metal3 s 59200 54620 60000 54860 6 io_oeb[36]
port 69 nsew signal output
rlabel metal3 s 59200 55436 60000 55676 6 io_oeb[37]
port 70 nsew signal output
rlabel metal3 s 59200 28236 60000 28476 6 io_oeb[3]
port 71 nsew signal output
rlabel metal3 s 59200 28916 60000 29156 6 io_oeb[4]
port 72 nsew signal output
rlabel metal3 s 59200 29732 60000 29972 6 io_oeb[5]
port 73 nsew signal output
rlabel metal3 s 59200 30548 60000 30788 6 io_oeb[6]
port 74 nsew signal output
rlabel metal3 s 59200 31364 60000 31604 6 io_oeb[7]
port 75 nsew signal output
rlabel metal3 s 59200 32180 60000 32420 6 io_oeb[8]
port 76 nsew signal output
rlabel metal3 s 59200 32996 60000 33236 6 io_oeb[9]
port 77 nsew signal output
rlabel metal2 s 31086 55200 31198 56000 6 io_out[0]
port 78 nsew signal output
rlabel metal2 s 38722 55200 38834 56000 6 io_out[10]
port 79 nsew signal output
rlabel metal2 s 39550 55200 39662 56000 6 io_out[11]
port 80 nsew signal output
rlabel metal2 s 40286 55200 40398 56000 6 io_out[12]
port 81 nsew signal output
rlabel metal2 s 41114 55200 41226 56000 6 io_out[13]
port 82 nsew signal output
rlabel metal2 s 41850 55200 41962 56000 6 io_out[14]
port 83 nsew signal output
rlabel metal2 s 42586 55200 42698 56000 6 io_out[15]
port 84 nsew signal output
rlabel metal2 s 43414 55200 43526 56000 6 io_out[16]
port 85 nsew signal output
rlabel metal2 s 44150 55200 44262 56000 6 io_out[17]
port 86 nsew signal output
rlabel metal2 s 44886 55200 44998 56000 6 io_out[18]
port 87 nsew signal output
rlabel metal2 s 45714 55200 45826 56000 6 io_out[19]
port 88 nsew signal output
rlabel metal2 s 31822 55200 31934 56000 6 io_out[1]
port 89 nsew signal output
rlabel metal2 s 46450 55200 46562 56000 6 io_out[20]
port 90 nsew signal output
rlabel metal2 s 47186 55200 47298 56000 6 io_out[21]
port 91 nsew signal output
rlabel metal2 s 48014 55200 48126 56000 6 io_out[22]
port 92 nsew signal output
rlabel metal2 s 48750 55200 48862 56000 6 io_out[23]
port 93 nsew signal output
rlabel metal2 s 49486 55200 49598 56000 6 io_out[24]
port 94 nsew signal output
rlabel metal2 s 50314 55200 50426 56000 6 io_out[25]
port 95 nsew signal output
rlabel metal2 s 51050 55200 51162 56000 6 io_out[26]
port 96 nsew signal output
rlabel metal2 s 51878 55200 51990 56000 6 io_out[27]
port 97 nsew signal output
rlabel metal2 s 52614 55200 52726 56000 6 io_out[28]
port 98 nsew signal output
rlabel metal2 s 53350 55200 53462 56000 6 io_out[29]
port 99 nsew signal output
rlabel metal2 s 32650 55200 32762 56000 6 io_out[2]
port 100 nsew signal output
rlabel metal2 s 54178 55200 54290 56000 6 io_out[30]
port 101 nsew signal output
rlabel metal2 s 54914 55200 55026 56000 6 io_out[31]
port 102 nsew signal output
rlabel metal2 s 55650 55200 55762 56000 6 io_out[32]
port 103 nsew signal output
rlabel metal2 s 56478 55200 56590 56000 6 io_out[33]
port 104 nsew signal output
rlabel metal2 s 57214 55200 57326 56000 6 io_out[34]
port 105 nsew signal output
rlabel metal2 s 57950 55200 58062 56000 6 io_out[35]
port 106 nsew signal output
rlabel metal2 s 58778 55200 58890 56000 6 io_out[36]
port 107 nsew signal output
rlabel metal2 s 59514 55200 59626 56000 6 io_out[37]
port 108 nsew signal output
rlabel metal2 s 33386 55200 33498 56000 6 io_out[3]
port 109 nsew signal output
rlabel metal2 s 34122 55200 34234 56000 6 io_out[4]
port 110 nsew signal output
rlabel metal2 s 34950 55200 35062 56000 6 io_out[5]
port 111 nsew signal output
rlabel metal2 s 35686 55200 35798 56000 6 io_out[6]
port 112 nsew signal output
rlabel metal2 s 36422 55200 36534 56000 6 io_out[7]
port 113 nsew signal output
rlabel metal2 s 37250 55200 37362 56000 6 io_out[8]
port 114 nsew signal output
rlabel metal2 s 37986 55200 38098 56000 6 io_out[9]
port 115 nsew signal output
rlabel metal3 s 0 356 800 596 6 la1_data_in[0]
port 116 nsew signal input
rlabel metal3 s 0 9060 800 9300 6 la1_data_in[10]
port 117 nsew signal input
rlabel metal3 s 0 9876 800 10116 6 la1_data_in[11]
port 118 nsew signal input
rlabel metal3 s 0 10828 800 11068 6 la1_data_in[12]
port 119 nsew signal input
rlabel metal3 s 0 11644 800 11884 6 la1_data_in[13]
port 120 nsew signal input
rlabel metal3 s 0 12596 800 12836 6 la1_data_in[14]
port 121 nsew signal input
rlabel metal3 s 0 13412 800 13652 6 la1_data_in[15]
port 122 nsew signal input
rlabel metal3 s 0 14364 800 14604 6 la1_data_in[16]
port 123 nsew signal input
rlabel metal3 s 0 15180 800 15420 6 la1_data_in[17]
port 124 nsew signal input
rlabel metal3 s 0 15996 800 16236 6 la1_data_in[18]
port 125 nsew signal input
rlabel metal3 s 0 16948 800 17188 6 la1_data_in[19]
port 126 nsew signal input
rlabel metal3 s 0 1172 800 1412 6 la1_data_in[1]
port 127 nsew signal input
rlabel metal3 s 0 17764 800 18004 6 la1_data_in[20]
port 128 nsew signal input
rlabel metal3 s 0 18716 800 18956 6 la1_data_in[21]
port 129 nsew signal input
rlabel metal3 s 0 19532 800 19772 6 la1_data_in[22]
port 130 nsew signal input
rlabel metal3 s 0 20484 800 20724 6 la1_data_in[23]
port 131 nsew signal input
rlabel metal3 s 0 21300 800 21540 6 la1_data_in[24]
port 132 nsew signal input
rlabel metal3 s 0 22116 800 22356 6 la1_data_in[25]
port 133 nsew signal input
rlabel metal3 s 0 23068 800 23308 6 la1_data_in[26]
port 134 nsew signal input
rlabel metal3 s 0 23884 800 24124 6 la1_data_in[27]
port 135 nsew signal input
rlabel metal3 s 0 24836 800 25076 6 la1_data_in[28]
port 136 nsew signal input
rlabel metal3 s 0 25652 800 25892 6 la1_data_in[29]
port 137 nsew signal input
rlabel metal3 s 0 1988 800 2228 6 la1_data_in[2]
port 138 nsew signal input
rlabel metal3 s 0 26604 800 26844 6 la1_data_in[30]
port 139 nsew signal input
rlabel metal3 s 0 27420 800 27660 6 la1_data_in[31]
port 140 nsew signal input
rlabel metal3 s 0 2940 800 3180 6 la1_data_in[3]
port 141 nsew signal input
rlabel metal3 s 0 3756 800 3996 6 la1_data_in[4]
port 142 nsew signal input
rlabel metal3 s 0 4708 800 4948 6 la1_data_in[5]
port 143 nsew signal input
rlabel metal3 s 0 5524 800 5764 6 la1_data_in[6]
port 144 nsew signal input
rlabel metal3 s 0 6476 800 6716 6 la1_data_in[7]
port 145 nsew signal input
rlabel metal3 s 0 7292 800 7532 6 la1_data_in[8]
port 146 nsew signal input
rlabel metal3 s 0 8108 800 8348 6 la1_data_in[9]
port 147 nsew signal input
rlabel metal3 s 0 28372 800 28612 6 la1_data_out[0]
port 148 nsew signal output
rlabel metal3 s 0 37076 800 37316 6 la1_data_out[10]
port 149 nsew signal output
rlabel metal3 s 0 37892 800 38132 6 la1_data_out[11]
port 150 nsew signal output
rlabel metal3 s 0 38844 800 39084 6 la1_data_out[12]
port 151 nsew signal output
rlabel metal3 s 0 39660 800 39900 6 la1_data_out[13]
port 152 nsew signal output
rlabel metal3 s 0 40612 800 40852 6 la1_data_out[14]
port 153 nsew signal output
rlabel metal3 s 0 41428 800 41668 6 la1_data_out[15]
port 154 nsew signal output
rlabel metal3 s 0 42380 800 42620 6 la1_data_out[16]
port 155 nsew signal output
rlabel metal3 s 0 43196 800 43436 6 la1_data_out[17]
port 156 nsew signal output
rlabel metal3 s 0 44012 800 44252 6 la1_data_out[18]
port 157 nsew signal output
rlabel metal3 s 0 44964 800 45204 6 la1_data_out[19]
port 158 nsew signal output
rlabel metal3 s 0 29188 800 29428 6 la1_data_out[1]
port 159 nsew signal output
rlabel metal3 s 0 45780 800 46020 6 la1_data_out[20]
port 160 nsew signal output
rlabel metal3 s 0 46732 800 46972 6 la1_data_out[21]
port 161 nsew signal output
rlabel metal3 s 0 47548 800 47788 6 la1_data_out[22]
port 162 nsew signal output
rlabel metal3 s 0 48500 800 48740 6 la1_data_out[23]
port 163 nsew signal output
rlabel metal3 s 0 49316 800 49556 6 la1_data_out[24]
port 164 nsew signal output
rlabel metal3 s 0 50132 800 50372 6 la1_data_out[25]
port 165 nsew signal output
rlabel metal3 s 0 51084 800 51324 6 la1_data_out[26]
port 166 nsew signal output
rlabel metal3 s 0 51900 800 52140 6 la1_data_out[27]
port 167 nsew signal output
rlabel metal3 s 0 52852 800 53092 6 la1_data_out[28]
port 168 nsew signal output
rlabel metal3 s 0 53668 800 53908 6 la1_data_out[29]
port 169 nsew signal output
rlabel metal3 s 0 30004 800 30244 6 la1_data_out[2]
port 170 nsew signal output
rlabel metal3 s 0 54620 800 54860 6 la1_data_out[30]
port 171 nsew signal output
rlabel metal3 s 0 55436 800 55676 6 la1_data_out[31]
port 172 nsew signal output
rlabel metal3 s 0 30956 800 31196 6 la1_data_out[3]
port 173 nsew signal output
rlabel metal3 s 0 31772 800 32012 6 la1_data_out[4]
port 174 nsew signal output
rlabel metal3 s 0 32724 800 32964 6 la1_data_out[5]
port 175 nsew signal output
rlabel metal3 s 0 33540 800 33780 6 la1_data_out[6]
port 176 nsew signal output
rlabel metal3 s 0 34492 800 34732 6 la1_data_out[7]
port 177 nsew signal output
rlabel metal3 s 0 35308 800 35548 6 la1_data_out[8]
port 178 nsew signal output
rlabel metal3 s 0 36124 800 36364 6 la1_data_out[9]
port 179 nsew signal output
rlabel metal3 s 59200 220 60000 460 6 la1_oenb[0]
port 180 nsew signal input
rlabel metal3 s 59200 8108 60000 8348 6 la1_oenb[10]
port 181 nsew signal input
rlabel metal3 s 59200 8924 60000 9164 6 la1_oenb[11]
port 182 nsew signal input
rlabel metal3 s 59200 9740 60000 9980 6 la1_oenb[12]
port 183 nsew signal input
rlabel metal3 s 59200 10556 60000 10796 6 la1_oenb[13]
port 184 nsew signal input
rlabel metal3 s 59200 11372 60000 11612 6 la1_oenb[14]
port 185 nsew signal input
rlabel metal3 s 59200 12188 60000 12428 6 la1_oenb[15]
port 186 nsew signal input
rlabel metal3 s 59200 13004 60000 13244 6 la1_oenb[16]
port 187 nsew signal input
rlabel metal3 s 59200 13820 60000 14060 6 la1_oenb[17]
port 188 nsew signal input
rlabel metal3 s 59200 14500 60000 14740 6 la1_oenb[18]
port 189 nsew signal input
rlabel metal3 s 59200 15316 60000 15556 6 la1_oenb[19]
port 190 nsew signal input
rlabel metal3 s 59200 900 60000 1140 6 la1_oenb[1]
port 191 nsew signal input
rlabel metal3 s 59200 16132 60000 16372 6 la1_oenb[20]
port 192 nsew signal input
rlabel metal3 s 59200 16948 60000 17188 6 la1_oenb[21]
port 193 nsew signal input
rlabel metal3 s 59200 17764 60000 18004 6 la1_oenb[22]
port 194 nsew signal input
rlabel metal3 s 59200 18580 60000 18820 6 la1_oenb[23]
port 195 nsew signal input
rlabel metal3 s 59200 19396 60000 19636 6 la1_oenb[24]
port 196 nsew signal input
rlabel metal3 s 59200 20212 60000 20452 6 la1_oenb[25]
port 197 nsew signal input
rlabel metal3 s 59200 21028 60000 21268 6 la1_oenb[26]
port 198 nsew signal input
rlabel metal3 s 59200 21708 60000 21948 6 la1_oenb[27]
port 199 nsew signal input
rlabel metal3 s 59200 22524 60000 22764 6 la1_oenb[28]
port 200 nsew signal input
rlabel metal3 s 59200 23340 60000 23580 6 la1_oenb[29]
port 201 nsew signal input
rlabel metal3 s 59200 1716 60000 1956 6 la1_oenb[2]
port 202 nsew signal input
rlabel metal3 s 59200 24156 60000 24396 6 la1_oenb[30]
port 203 nsew signal input
rlabel metal3 s 59200 24972 60000 25212 6 la1_oenb[31]
port 204 nsew signal input
rlabel metal3 s 59200 2532 60000 2772 6 la1_oenb[3]
port 205 nsew signal input
rlabel metal3 s 59200 3348 60000 3588 6 la1_oenb[4]
port 206 nsew signal input
rlabel metal3 s 59200 4164 60000 4404 6 la1_oenb[5]
port 207 nsew signal input
rlabel metal3 s 59200 4980 60000 5220 6 la1_oenb[6]
port 208 nsew signal input
rlabel metal3 s 59200 5796 60000 6036 6 la1_oenb[7]
port 209 nsew signal input
rlabel metal3 s 59200 6612 60000 6852 6 la1_oenb[8]
port 210 nsew signal input
rlabel metal3 s 59200 7292 60000 7532 6 la1_oenb[9]
port 211 nsew signal input
rlabel metal4 s 4208 496 4528 53360 6 vccd1
port 212 nsew power input
rlabel metal4 s 34928 496 35248 53360 6 vccd1
port 212 nsew power input
rlabel metal4 s 19568 496 19888 53360 6 vssd1
port 213 nsew ground input
rlabel metal4 s 50288 496 50608 53360 6 vssd1
port 213 nsew ground input
rlabel metal2 s 1094 55200 1206 56000 6 wb_clk_i
port 214 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 60000 56000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 12996724
string GDS_FILE /openlane/designs/wrapped_vgademo_on_fpga/runs/RUN_2022.03.20_01.02.09/results/finishing/wrapped_vgademo_on_fpga.magic.gds
string GDS_START 1050072
<< end >>

