magic
tech sky130A
magscale 1 2
timestamp 1647761360
<< obsli1 >>
rect 1104 527 58880 57681
<< obsm1 >>
rect 566 212 59326 58064
<< metal2 >>
rect 542 59200 654 60000
rect 1738 59200 1850 60000
rect 2934 59200 3046 60000
rect 4130 59200 4242 60000
rect 5418 59200 5530 60000
rect 6614 59200 6726 60000
rect 7810 59200 7922 60000
rect 9098 59200 9210 60000
rect 10294 59200 10406 60000
rect 11490 59200 11602 60000
rect 12778 59200 12890 60000
rect 13974 59200 14086 60000
rect 15170 59200 15282 60000
rect 16366 59200 16478 60000
rect 17654 59200 17766 60000
rect 18850 59200 18962 60000
rect 20046 59200 20158 60000
rect 21334 59200 21446 60000
rect 22530 59200 22642 60000
rect 23726 59200 23838 60000
rect 25014 59200 25126 60000
rect 26210 59200 26322 60000
rect 27406 59200 27518 60000
rect 28694 59200 28806 60000
rect 29890 59200 30002 60000
rect 31086 59200 31198 60000
rect 32282 59200 32394 60000
rect 33570 59200 33682 60000
rect 34766 59200 34878 60000
rect 35962 59200 36074 60000
rect 37250 59200 37362 60000
rect 38446 59200 38558 60000
rect 39642 59200 39754 60000
rect 40930 59200 41042 60000
rect 42126 59200 42238 60000
rect 43322 59200 43434 60000
rect 44610 59200 44722 60000
rect 45806 59200 45918 60000
rect 47002 59200 47114 60000
rect 48198 59200 48310 60000
rect 49486 59200 49598 60000
rect 50682 59200 50794 60000
rect 51878 59200 51990 60000
rect 53166 59200 53278 60000
rect 54362 59200 54474 60000
rect 55558 59200 55670 60000
rect 56846 59200 56958 60000
rect 58042 59200 58154 60000
rect 59238 59200 59350 60000
rect 3302 0 3414 800
rect 9926 0 10038 800
rect 16550 0 16662 800
rect 23266 0 23378 800
rect 29890 0 30002 800
rect 36606 0 36718 800
rect 43230 0 43342 800
rect 49946 0 50058 800
rect 56570 0 56682 800
<< obsm2 >>
rect 710 59144 1682 59537
rect 1906 59144 2878 59537
rect 3102 59144 4074 59537
rect 4298 59144 5362 59537
rect 5586 59144 6558 59537
rect 6782 59144 7754 59537
rect 7978 59144 9042 59537
rect 9266 59144 10238 59537
rect 10462 59144 11434 59537
rect 11658 59144 12722 59537
rect 12946 59144 13918 59537
rect 14142 59144 15114 59537
rect 15338 59144 16310 59537
rect 16534 59144 17598 59537
rect 17822 59144 18794 59537
rect 19018 59144 19990 59537
rect 20214 59144 21278 59537
rect 21502 59144 22474 59537
rect 22698 59144 23670 59537
rect 23894 59144 24958 59537
rect 25182 59144 26154 59537
rect 26378 59144 27350 59537
rect 27574 59144 28638 59537
rect 28862 59144 29834 59537
rect 30058 59144 31030 59537
rect 31254 59144 32226 59537
rect 32450 59144 33514 59537
rect 33738 59144 34710 59537
rect 34934 59144 35906 59537
rect 36130 59144 37194 59537
rect 37418 59144 38390 59537
rect 38614 59144 39586 59537
rect 39810 59144 40874 59537
rect 41098 59144 42070 59537
rect 42294 59144 43266 59537
rect 43490 59144 44554 59537
rect 44778 59144 45750 59537
rect 45974 59144 46946 59537
rect 47170 59144 48142 59537
rect 48366 59144 49430 59537
rect 49654 59144 50626 59537
rect 50850 59144 51822 59537
rect 52046 59144 53110 59537
rect 53334 59144 54306 59537
rect 54530 59144 55502 59537
rect 55726 59144 56790 59537
rect 57014 59144 57986 59537
rect 58210 59144 59182 59537
rect 572 856 59320 59144
rect 572 206 3246 856
rect 3470 206 9870 856
rect 10094 206 16494 856
rect 16718 206 23210 856
rect 23434 206 29834 856
rect 30058 206 36550 856
rect 36774 206 43174 856
rect 43398 206 49890 856
rect 50114 206 56514 856
rect 56738 206 59320 856
<< metal3 >>
rect 0 59380 800 59620
rect 59200 59380 60000 59620
rect 0 58564 800 58804
rect 59200 58700 60000 58940
rect 0 57748 800 57988
rect 59200 57884 60000 58124
rect 0 56932 800 57172
rect 59200 57204 60000 57444
rect 0 56116 800 56356
rect 59200 56388 60000 56628
rect 59200 55708 60000 55948
rect 0 55300 800 55540
rect 59200 54892 60000 55132
rect 0 54484 800 54724
rect 59200 54212 60000 54452
rect 0 53668 800 53908
rect 59200 53532 60000 53772
rect 0 52852 800 53092
rect 59200 52716 60000 52956
rect 0 52036 800 52276
rect 59200 52036 60000 52276
rect 0 51220 800 51460
rect 59200 51220 60000 51460
rect 0 50404 800 50644
rect 59200 50540 60000 50780
rect 0 49588 800 49828
rect 59200 49724 60000 49964
rect 0 48772 800 49012
rect 59200 49044 60000 49284
rect 0 47956 800 48196
rect 59200 48228 60000 48468
rect 59200 47548 60000 47788
rect 0 47140 800 47380
rect 59200 46868 60000 47108
rect 0 46324 800 46564
rect 59200 46052 60000 46292
rect 0 45508 800 45748
rect 59200 45372 60000 45612
rect 0 44692 800 44932
rect 59200 44556 60000 44796
rect 0 43876 800 44116
rect 59200 43876 60000 44116
rect 0 43060 800 43300
rect 59200 43060 60000 43300
rect 0 42244 800 42484
rect 59200 42380 60000 42620
rect 0 41428 800 41668
rect 59200 41564 60000 41804
rect 0 40612 800 40852
rect 59200 40884 60000 41124
rect 59200 40204 60000 40444
rect 0 39660 800 39900
rect 59200 39388 60000 39628
rect 0 38844 800 39084
rect 59200 38708 60000 38948
rect 0 38028 800 38268
rect 59200 37892 60000 38132
rect 0 37212 800 37452
rect 59200 37212 60000 37452
rect 0 36396 800 36636
rect 59200 36396 60000 36636
rect 0 35580 800 35820
rect 59200 35716 60000 35956
rect 0 34764 800 35004
rect 59200 34900 60000 35140
rect 0 33948 800 34188
rect 59200 34220 60000 34460
rect 59200 33540 60000 33780
rect 0 33132 800 33372
rect 59200 32724 60000 32964
rect 0 32316 800 32556
rect 59200 32044 60000 32284
rect 0 31500 800 31740
rect 59200 31228 60000 31468
rect 0 30684 800 30924
rect 59200 30548 60000 30788
rect 0 29868 800 30108
rect 59200 29732 60000 29972
rect 0 29052 800 29292
rect 59200 29052 60000 29292
rect 0 28236 800 28476
rect 59200 28236 60000 28476
rect 0 27420 800 27660
rect 59200 27556 60000 27796
rect 0 26604 800 26844
rect 59200 26876 60000 27116
rect 0 25788 800 26028
rect 59200 26060 60000 26300
rect 59200 25380 60000 25620
rect 0 24972 800 25212
rect 59200 24564 60000 24804
rect 0 24156 800 24396
rect 59200 23884 60000 24124
rect 0 23340 800 23580
rect 59200 23068 60000 23308
rect 0 22524 800 22764
rect 59200 22388 60000 22628
rect 0 21708 800 21948
rect 59200 21572 60000 21812
rect 0 20892 800 21132
rect 59200 20892 60000 21132
rect 0 19940 800 20180
rect 59200 20212 60000 20452
rect 0 19124 800 19364
rect 59200 19396 60000 19636
rect 59200 18716 60000 18956
rect 0 18308 800 18548
rect 59200 17900 60000 18140
rect 0 17492 800 17732
rect 59200 17220 60000 17460
rect 0 16676 800 16916
rect 59200 16404 60000 16644
rect 0 15860 800 16100
rect 59200 15724 60000 15964
rect 0 15044 800 15284
rect 59200 14908 60000 15148
rect 0 14228 800 14468
rect 59200 14228 60000 14468
rect 0 13412 800 13652
rect 59200 13548 60000 13788
rect 0 12596 800 12836
rect 59200 12732 60000 12972
rect 0 11780 800 12020
rect 59200 12052 60000 12292
rect 0 10964 800 11204
rect 59200 11236 60000 11476
rect 59200 10556 60000 10796
rect 0 10148 800 10388
rect 59200 9740 60000 9980
rect 0 9332 800 9572
rect 59200 9060 60000 9300
rect 0 8516 800 8756
rect 59200 8244 60000 8484
rect 0 7700 800 7940
rect 59200 7564 60000 7804
rect 0 6884 800 7124
rect 59200 6884 60000 7124
rect 0 6068 800 6308
rect 59200 6068 60000 6308
rect 0 5252 800 5492
rect 59200 5388 60000 5628
rect 0 4436 800 4676
rect 59200 4572 60000 4812
rect 0 3620 800 3860
rect 59200 3892 60000 4132
rect 0 2804 800 3044
rect 59200 3076 60000 3316
rect 59200 2396 60000 2636
rect 0 1988 800 2228
rect 59200 1580 60000 1820
rect 0 1172 800 1412
rect 59200 900 60000 1140
rect 0 356 800 596
rect 59200 220 60000 460
<< obsm3 >>
rect 880 59300 59120 59533
rect 800 59020 59200 59300
rect 800 58884 59120 59020
rect 880 58620 59120 58884
rect 880 58484 59200 58620
rect 800 58204 59200 58484
rect 800 58068 59120 58204
rect 880 57804 59120 58068
rect 880 57668 59200 57804
rect 800 57524 59200 57668
rect 800 57252 59120 57524
rect 880 57124 59120 57252
rect 880 56852 59200 57124
rect 800 56708 59200 56852
rect 800 56436 59120 56708
rect 880 56308 59120 56436
rect 880 56036 59200 56308
rect 800 56028 59200 56036
rect 800 55628 59120 56028
rect 800 55620 59200 55628
rect 880 55220 59200 55620
rect 800 55212 59200 55220
rect 800 54812 59120 55212
rect 800 54804 59200 54812
rect 880 54532 59200 54804
rect 880 54404 59120 54532
rect 800 54132 59120 54404
rect 800 53988 59200 54132
rect 880 53852 59200 53988
rect 880 53588 59120 53852
rect 800 53452 59120 53588
rect 800 53172 59200 53452
rect 880 53036 59200 53172
rect 880 52772 59120 53036
rect 800 52636 59120 52772
rect 800 52356 59200 52636
rect 880 51956 59120 52356
rect 800 51540 59200 51956
rect 880 51140 59120 51540
rect 800 50860 59200 51140
rect 800 50724 59120 50860
rect 880 50460 59120 50724
rect 880 50324 59200 50460
rect 800 50044 59200 50324
rect 800 49908 59120 50044
rect 880 49644 59120 49908
rect 880 49508 59200 49644
rect 800 49364 59200 49508
rect 800 49092 59120 49364
rect 880 48964 59120 49092
rect 880 48692 59200 48964
rect 800 48548 59200 48692
rect 800 48276 59120 48548
rect 880 48148 59120 48276
rect 880 47876 59200 48148
rect 800 47868 59200 47876
rect 800 47468 59120 47868
rect 800 47460 59200 47468
rect 880 47188 59200 47460
rect 880 47060 59120 47188
rect 800 46788 59120 47060
rect 800 46644 59200 46788
rect 880 46372 59200 46644
rect 880 46244 59120 46372
rect 800 45972 59120 46244
rect 800 45828 59200 45972
rect 880 45692 59200 45828
rect 880 45428 59120 45692
rect 800 45292 59120 45428
rect 800 45012 59200 45292
rect 880 44876 59200 45012
rect 880 44612 59120 44876
rect 800 44476 59120 44612
rect 800 44196 59200 44476
rect 880 43796 59120 44196
rect 800 43380 59200 43796
rect 880 42980 59120 43380
rect 800 42700 59200 42980
rect 800 42564 59120 42700
rect 880 42300 59120 42564
rect 880 42164 59200 42300
rect 800 41884 59200 42164
rect 800 41748 59120 41884
rect 880 41484 59120 41748
rect 880 41348 59200 41484
rect 800 41204 59200 41348
rect 800 40932 59120 41204
rect 880 40804 59120 40932
rect 880 40532 59200 40804
rect 800 40524 59200 40532
rect 800 40124 59120 40524
rect 800 39980 59200 40124
rect 880 39708 59200 39980
rect 880 39580 59120 39708
rect 800 39308 59120 39580
rect 800 39164 59200 39308
rect 880 39028 59200 39164
rect 880 38764 59120 39028
rect 800 38628 59120 38764
rect 800 38348 59200 38628
rect 880 38212 59200 38348
rect 880 37948 59120 38212
rect 800 37812 59120 37948
rect 800 37532 59200 37812
rect 880 37132 59120 37532
rect 800 36716 59200 37132
rect 880 36316 59120 36716
rect 800 36036 59200 36316
rect 800 35900 59120 36036
rect 880 35636 59120 35900
rect 880 35500 59200 35636
rect 800 35220 59200 35500
rect 800 35084 59120 35220
rect 880 34820 59120 35084
rect 880 34684 59200 34820
rect 800 34540 59200 34684
rect 800 34268 59120 34540
rect 880 34140 59120 34268
rect 880 33868 59200 34140
rect 800 33860 59200 33868
rect 800 33460 59120 33860
rect 800 33452 59200 33460
rect 880 33052 59200 33452
rect 800 33044 59200 33052
rect 800 32644 59120 33044
rect 800 32636 59200 32644
rect 880 32364 59200 32636
rect 880 32236 59120 32364
rect 800 31964 59120 32236
rect 800 31820 59200 31964
rect 880 31548 59200 31820
rect 880 31420 59120 31548
rect 800 31148 59120 31420
rect 800 31004 59200 31148
rect 880 30868 59200 31004
rect 880 30604 59120 30868
rect 800 30468 59120 30604
rect 800 30188 59200 30468
rect 880 30052 59200 30188
rect 880 29788 59120 30052
rect 800 29652 59120 29788
rect 800 29372 59200 29652
rect 880 28972 59120 29372
rect 800 28556 59200 28972
rect 880 28156 59120 28556
rect 800 27876 59200 28156
rect 800 27740 59120 27876
rect 880 27476 59120 27740
rect 880 27340 59200 27476
rect 800 27196 59200 27340
rect 800 26924 59120 27196
rect 880 26796 59120 26924
rect 880 26524 59200 26796
rect 800 26380 59200 26524
rect 800 26108 59120 26380
rect 880 25980 59120 26108
rect 880 25708 59200 25980
rect 800 25700 59200 25708
rect 800 25300 59120 25700
rect 800 25292 59200 25300
rect 880 24892 59200 25292
rect 800 24884 59200 24892
rect 800 24484 59120 24884
rect 800 24476 59200 24484
rect 880 24204 59200 24476
rect 880 24076 59120 24204
rect 800 23804 59120 24076
rect 800 23660 59200 23804
rect 880 23388 59200 23660
rect 880 23260 59120 23388
rect 800 22988 59120 23260
rect 800 22844 59200 22988
rect 880 22708 59200 22844
rect 880 22444 59120 22708
rect 800 22308 59120 22444
rect 800 22028 59200 22308
rect 880 21892 59200 22028
rect 880 21628 59120 21892
rect 800 21492 59120 21628
rect 800 21212 59200 21492
rect 880 20812 59120 21212
rect 800 20532 59200 20812
rect 800 20260 59120 20532
rect 880 20132 59120 20260
rect 880 19860 59200 20132
rect 800 19716 59200 19860
rect 800 19444 59120 19716
rect 880 19316 59120 19444
rect 880 19044 59200 19316
rect 800 19036 59200 19044
rect 800 18636 59120 19036
rect 800 18628 59200 18636
rect 880 18228 59200 18628
rect 800 18220 59200 18228
rect 800 17820 59120 18220
rect 800 17812 59200 17820
rect 880 17540 59200 17812
rect 880 17412 59120 17540
rect 800 17140 59120 17412
rect 800 16996 59200 17140
rect 880 16724 59200 16996
rect 880 16596 59120 16724
rect 800 16324 59120 16596
rect 800 16180 59200 16324
rect 880 16044 59200 16180
rect 880 15780 59120 16044
rect 800 15644 59120 15780
rect 800 15364 59200 15644
rect 880 15228 59200 15364
rect 880 14964 59120 15228
rect 800 14828 59120 14964
rect 800 14548 59200 14828
rect 880 14148 59120 14548
rect 800 13868 59200 14148
rect 800 13732 59120 13868
rect 880 13468 59120 13732
rect 880 13332 59200 13468
rect 800 13052 59200 13332
rect 800 12916 59120 13052
rect 880 12652 59120 12916
rect 880 12516 59200 12652
rect 800 12372 59200 12516
rect 800 12100 59120 12372
rect 880 11972 59120 12100
rect 880 11700 59200 11972
rect 800 11556 59200 11700
rect 800 11284 59120 11556
rect 880 11156 59120 11284
rect 880 10884 59200 11156
rect 800 10876 59200 10884
rect 800 10476 59120 10876
rect 800 10468 59200 10476
rect 880 10068 59200 10468
rect 800 10060 59200 10068
rect 800 9660 59120 10060
rect 800 9652 59200 9660
rect 880 9380 59200 9652
rect 880 9252 59120 9380
rect 800 8980 59120 9252
rect 800 8836 59200 8980
rect 880 8564 59200 8836
rect 880 8436 59120 8564
rect 800 8164 59120 8436
rect 800 8020 59200 8164
rect 880 7884 59200 8020
rect 880 7620 59120 7884
rect 800 7484 59120 7620
rect 800 7204 59200 7484
rect 880 6804 59120 7204
rect 800 6388 59200 6804
rect 880 5988 59120 6388
rect 800 5708 59200 5988
rect 800 5572 59120 5708
rect 880 5308 59120 5572
rect 880 5172 59200 5308
rect 800 4892 59200 5172
rect 800 4756 59120 4892
rect 880 4492 59120 4756
rect 880 4356 59200 4492
rect 800 4212 59200 4356
rect 800 3940 59120 4212
rect 880 3812 59120 3940
rect 880 3540 59200 3812
rect 800 3396 59200 3540
rect 800 3124 59120 3396
rect 880 2996 59120 3124
rect 880 2724 59200 2996
rect 800 2716 59200 2724
rect 800 2316 59120 2716
rect 800 2308 59200 2316
rect 880 1908 59200 2308
rect 800 1900 59200 1908
rect 800 1500 59120 1900
rect 800 1492 59200 1500
rect 880 1220 59200 1492
rect 880 1092 59120 1220
rect 800 820 59120 1092
rect 800 676 59200 820
rect 880 540 59200 676
rect 880 511 59120 540
<< metal4 >>
rect 4208 496 4528 57712
rect 19568 496 19888 57712
rect 34928 496 35248 57712
rect 50288 496 50608 57712
<< obsm4 >>
rect 4659 1395 19488 52597
rect 19968 1395 34848 52597
rect 35328 1395 48517 52597
<< labels >>
rlabel metal2 s 542 59200 654 60000 6 active
port 1 nsew signal input
rlabel metal2 s 2934 59200 3046 60000 6 io_in[0]
port 2 nsew signal input
rlabel metal2 s 15170 59200 15282 60000 6 io_in[10]
port 3 nsew signal input
rlabel metal2 s 16366 59200 16478 60000 6 io_in[11]
port 4 nsew signal input
rlabel metal2 s 17654 59200 17766 60000 6 io_in[12]
port 5 nsew signal input
rlabel metal2 s 18850 59200 18962 60000 6 io_in[13]
port 6 nsew signal input
rlabel metal2 s 20046 59200 20158 60000 6 io_in[14]
port 7 nsew signal input
rlabel metal2 s 21334 59200 21446 60000 6 io_in[15]
port 8 nsew signal input
rlabel metal2 s 22530 59200 22642 60000 6 io_in[16]
port 9 nsew signal input
rlabel metal2 s 23726 59200 23838 60000 6 io_in[17]
port 10 nsew signal input
rlabel metal2 s 25014 59200 25126 60000 6 io_in[18]
port 11 nsew signal input
rlabel metal2 s 26210 59200 26322 60000 6 io_in[19]
port 12 nsew signal input
rlabel metal2 s 4130 59200 4242 60000 6 io_in[1]
port 13 nsew signal input
rlabel metal2 s 27406 59200 27518 60000 6 io_in[20]
port 14 nsew signal input
rlabel metal2 s 28694 59200 28806 60000 6 io_in[21]
port 15 nsew signal input
rlabel metal2 s 29890 59200 30002 60000 6 io_in[22]
port 16 nsew signal input
rlabel metal2 s 31086 59200 31198 60000 6 io_in[23]
port 17 nsew signal input
rlabel metal2 s 32282 59200 32394 60000 6 io_in[24]
port 18 nsew signal input
rlabel metal2 s 33570 59200 33682 60000 6 io_in[25]
port 19 nsew signal input
rlabel metal2 s 34766 59200 34878 60000 6 io_in[26]
port 20 nsew signal input
rlabel metal2 s 35962 59200 36074 60000 6 io_in[27]
port 21 nsew signal input
rlabel metal2 s 37250 59200 37362 60000 6 io_in[28]
port 22 nsew signal input
rlabel metal2 s 38446 59200 38558 60000 6 io_in[29]
port 23 nsew signal input
rlabel metal2 s 5418 59200 5530 60000 6 io_in[2]
port 24 nsew signal input
rlabel metal2 s 39642 59200 39754 60000 6 io_in[30]
port 25 nsew signal input
rlabel metal2 s 40930 59200 41042 60000 6 io_in[31]
port 26 nsew signal input
rlabel metal2 s 42126 59200 42238 60000 6 io_in[32]
port 27 nsew signal input
rlabel metal2 s 43322 59200 43434 60000 6 io_in[33]
port 28 nsew signal input
rlabel metal2 s 44610 59200 44722 60000 6 io_in[34]
port 29 nsew signal input
rlabel metal2 s 45806 59200 45918 60000 6 io_in[35]
port 30 nsew signal input
rlabel metal2 s 47002 59200 47114 60000 6 io_in[36]
port 31 nsew signal input
rlabel metal2 s 48198 59200 48310 60000 6 io_in[37]
port 32 nsew signal input
rlabel metal2 s 6614 59200 6726 60000 6 io_in[3]
port 33 nsew signal input
rlabel metal2 s 7810 59200 7922 60000 6 io_in[4]
port 34 nsew signal input
rlabel metal2 s 9098 59200 9210 60000 6 io_in[5]
port 35 nsew signal input
rlabel metal2 s 10294 59200 10406 60000 6 io_in[6]
port 36 nsew signal input
rlabel metal2 s 11490 59200 11602 60000 6 io_in[7]
port 37 nsew signal input
rlabel metal2 s 12778 59200 12890 60000 6 io_in[8]
port 38 nsew signal input
rlabel metal2 s 13974 59200 14086 60000 6 io_in[9]
port 39 nsew signal input
rlabel metal3 s 59200 23884 60000 24124 6 io_oeb[0]
port 40 nsew signal output
rlabel metal3 s 59200 31228 60000 31468 6 io_oeb[10]
port 41 nsew signal output
rlabel metal3 s 59200 32044 60000 32284 6 io_oeb[11]
port 42 nsew signal output
rlabel metal3 s 59200 32724 60000 32964 6 io_oeb[12]
port 43 nsew signal output
rlabel metal3 s 59200 33540 60000 33780 6 io_oeb[13]
port 44 nsew signal output
rlabel metal3 s 59200 34220 60000 34460 6 io_oeb[14]
port 45 nsew signal output
rlabel metal3 s 59200 34900 60000 35140 6 io_oeb[15]
port 46 nsew signal output
rlabel metal3 s 59200 35716 60000 35956 6 io_oeb[16]
port 47 nsew signal output
rlabel metal3 s 59200 36396 60000 36636 6 io_oeb[17]
port 48 nsew signal output
rlabel metal3 s 59200 37212 60000 37452 6 io_oeb[18]
port 49 nsew signal output
rlabel metal3 s 59200 37892 60000 38132 6 io_oeb[19]
port 50 nsew signal output
rlabel metal3 s 59200 24564 60000 24804 6 io_oeb[1]
port 51 nsew signal output
rlabel metal3 s 59200 38708 60000 38948 6 io_oeb[20]
port 52 nsew signal output
rlabel metal3 s 59200 39388 60000 39628 6 io_oeb[21]
port 53 nsew signal output
rlabel metal3 s 59200 40204 60000 40444 6 io_oeb[22]
port 54 nsew signal output
rlabel metal3 s 59200 40884 60000 41124 6 io_oeb[23]
port 55 nsew signal output
rlabel metal3 s 59200 41564 60000 41804 6 io_oeb[24]
port 56 nsew signal output
rlabel metal3 s 59200 42380 60000 42620 6 io_oeb[25]
port 57 nsew signal output
rlabel metal3 s 59200 43060 60000 43300 6 io_oeb[26]
port 58 nsew signal output
rlabel metal3 s 59200 43876 60000 44116 6 io_oeb[27]
port 59 nsew signal output
rlabel metal3 s 59200 44556 60000 44796 6 io_oeb[28]
port 60 nsew signal output
rlabel metal3 s 59200 45372 60000 45612 6 io_oeb[29]
port 61 nsew signal output
rlabel metal3 s 59200 25380 60000 25620 6 io_oeb[2]
port 62 nsew signal output
rlabel metal3 s 59200 46052 60000 46292 6 io_oeb[30]
port 63 nsew signal output
rlabel metal3 s 59200 46868 60000 47108 6 io_oeb[31]
port 64 nsew signal output
rlabel metal3 s 59200 47548 60000 47788 6 io_oeb[32]
port 65 nsew signal output
rlabel metal3 s 59200 48228 60000 48468 6 io_oeb[33]
port 66 nsew signal output
rlabel metal3 s 59200 49044 60000 49284 6 io_oeb[34]
port 67 nsew signal output
rlabel metal3 s 59200 49724 60000 49964 6 io_oeb[35]
port 68 nsew signal output
rlabel metal3 s 59200 50540 60000 50780 6 io_oeb[36]
port 69 nsew signal output
rlabel metal3 s 59200 51220 60000 51460 6 io_oeb[37]
port 70 nsew signal output
rlabel metal3 s 59200 26060 60000 26300 6 io_oeb[3]
port 71 nsew signal output
rlabel metal3 s 59200 26876 60000 27116 6 io_oeb[4]
port 72 nsew signal output
rlabel metal3 s 59200 27556 60000 27796 6 io_oeb[5]
port 73 nsew signal output
rlabel metal3 s 59200 28236 60000 28476 6 io_oeb[6]
port 74 nsew signal output
rlabel metal3 s 59200 29052 60000 29292 6 io_oeb[7]
port 75 nsew signal output
rlabel metal3 s 59200 29732 60000 29972 6 io_oeb[8]
port 76 nsew signal output
rlabel metal3 s 59200 30548 60000 30788 6 io_oeb[9]
port 77 nsew signal output
rlabel metal2 s 3302 0 3414 800 6 io_out[0]
port 78 nsew signal output
rlabel metal2 s 49486 59200 49598 60000 6 io_out[10]
port 79 nsew signal output
rlabel metal3 s 59200 54212 60000 54452 6 io_out[11]
port 80 nsew signal output
rlabel metal3 s 59200 54892 60000 55132 6 io_out[12]
port 81 nsew signal output
rlabel metal2 s 29890 0 30002 800 6 io_out[13]
port 82 nsew signal output
rlabel metal2 s 36606 0 36718 800 6 io_out[14]
port 83 nsew signal output
rlabel metal2 s 50682 59200 50794 60000 6 io_out[15]
port 84 nsew signal output
rlabel metal3 s 59200 55708 60000 55948 6 io_out[16]
port 85 nsew signal output
rlabel metal3 s 59200 56388 60000 56628 6 io_out[17]
port 86 nsew signal output
rlabel metal3 s 59200 57204 60000 57444 6 io_out[18]
port 87 nsew signal output
rlabel metal3 s 0 55300 800 55540 6 io_out[19]
port 88 nsew signal output
rlabel metal3 s 59200 52036 60000 52276 6 io_out[1]
port 89 nsew signal output
rlabel metal2 s 43230 0 43342 800 6 io_out[20]
port 90 nsew signal output
rlabel metal3 s 59200 57884 60000 58124 6 io_out[21]
port 91 nsew signal output
rlabel metal2 s 49946 0 50058 800 6 io_out[22]
port 92 nsew signal output
rlabel metal3 s 0 56116 800 56356 6 io_out[23]
port 93 nsew signal output
rlabel metal3 s 59200 58700 60000 58940 6 io_out[24]
port 94 nsew signal output
rlabel metal3 s 0 56932 800 57172 6 io_out[25]
port 95 nsew signal output
rlabel metal2 s 51878 59200 51990 60000 6 io_out[26]
port 96 nsew signal output
rlabel metal3 s 0 57748 800 57988 6 io_out[27]
port 97 nsew signal output
rlabel metal2 s 53166 59200 53278 60000 6 io_out[28]
port 98 nsew signal output
rlabel metal3 s 59200 59380 60000 59620 6 io_out[29]
port 99 nsew signal output
rlabel metal2 s 9926 0 10038 800 6 io_out[2]
port 100 nsew signal output
rlabel metal3 s 0 58564 800 58804 6 io_out[30]
port 101 nsew signal output
rlabel metal2 s 54362 59200 54474 60000 6 io_out[31]
port 102 nsew signal output
rlabel metal2 s 55558 59200 55670 60000 6 io_out[32]
port 103 nsew signal output
rlabel metal2 s 56846 59200 56958 60000 6 io_out[33]
port 104 nsew signal output
rlabel metal2 s 56570 0 56682 800 6 io_out[34]
port 105 nsew signal output
rlabel metal3 s 0 59380 800 59620 6 io_out[35]
port 106 nsew signal output
rlabel metal2 s 58042 59200 58154 60000 6 io_out[36]
port 107 nsew signal output
rlabel metal2 s 59238 59200 59350 60000 6 io_out[37]
port 108 nsew signal output
rlabel metal2 s 16550 0 16662 800 6 io_out[3]
port 109 nsew signal output
rlabel metal3 s 59200 52716 60000 52956 6 io_out[4]
port 110 nsew signal output
rlabel metal2 s 23266 0 23378 800 6 io_out[5]
port 111 nsew signal output
rlabel metal3 s 59200 53532 60000 53772 6 io_out[6]
port 112 nsew signal output
rlabel metal3 s 0 52852 800 53092 6 io_out[7]
port 113 nsew signal output
rlabel metal3 s 0 53668 800 53908 6 io_out[8]
port 114 nsew signal output
rlabel metal3 s 0 54484 800 54724 6 io_out[9]
port 115 nsew signal output
rlabel metal3 s 0 356 800 596 6 la1_data_in[0]
port 116 nsew signal input
rlabel metal3 s 0 8516 800 8756 6 la1_data_in[10]
port 117 nsew signal input
rlabel metal3 s 0 9332 800 9572 6 la1_data_in[11]
port 118 nsew signal input
rlabel metal3 s 0 10148 800 10388 6 la1_data_in[12]
port 119 nsew signal input
rlabel metal3 s 0 10964 800 11204 6 la1_data_in[13]
port 120 nsew signal input
rlabel metal3 s 0 11780 800 12020 6 la1_data_in[14]
port 121 nsew signal input
rlabel metal3 s 0 12596 800 12836 6 la1_data_in[15]
port 122 nsew signal input
rlabel metal3 s 0 13412 800 13652 6 la1_data_in[16]
port 123 nsew signal input
rlabel metal3 s 0 14228 800 14468 6 la1_data_in[17]
port 124 nsew signal input
rlabel metal3 s 0 15044 800 15284 6 la1_data_in[18]
port 125 nsew signal input
rlabel metal3 s 0 15860 800 16100 6 la1_data_in[19]
port 126 nsew signal input
rlabel metal3 s 0 1172 800 1412 6 la1_data_in[1]
port 127 nsew signal input
rlabel metal3 s 0 16676 800 16916 6 la1_data_in[20]
port 128 nsew signal input
rlabel metal3 s 0 17492 800 17732 6 la1_data_in[21]
port 129 nsew signal input
rlabel metal3 s 0 18308 800 18548 6 la1_data_in[22]
port 130 nsew signal input
rlabel metal3 s 0 19124 800 19364 6 la1_data_in[23]
port 131 nsew signal input
rlabel metal3 s 0 19940 800 20180 6 la1_data_in[24]
port 132 nsew signal input
rlabel metal3 s 0 20892 800 21132 6 la1_data_in[25]
port 133 nsew signal input
rlabel metal3 s 0 21708 800 21948 6 la1_data_in[26]
port 134 nsew signal input
rlabel metal3 s 0 22524 800 22764 6 la1_data_in[27]
port 135 nsew signal input
rlabel metal3 s 0 23340 800 23580 6 la1_data_in[28]
port 136 nsew signal input
rlabel metal3 s 0 24156 800 24396 6 la1_data_in[29]
port 137 nsew signal input
rlabel metal3 s 0 1988 800 2228 6 la1_data_in[2]
port 138 nsew signal input
rlabel metal3 s 0 24972 800 25212 6 la1_data_in[30]
port 139 nsew signal input
rlabel metal3 s 0 25788 800 26028 6 la1_data_in[31]
port 140 nsew signal input
rlabel metal3 s 0 2804 800 3044 6 la1_data_in[3]
port 141 nsew signal input
rlabel metal3 s 0 3620 800 3860 6 la1_data_in[4]
port 142 nsew signal input
rlabel metal3 s 0 4436 800 4676 6 la1_data_in[5]
port 143 nsew signal input
rlabel metal3 s 0 5252 800 5492 6 la1_data_in[6]
port 144 nsew signal input
rlabel metal3 s 0 6068 800 6308 6 la1_data_in[7]
port 145 nsew signal input
rlabel metal3 s 0 6884 800 7124 6 la1_data_in[8]
port 146 nsew signal input
rlabel metal3 s 0 7700 800 7940 6 la1_data_in[9]
port 147 nsew signal input
rlabel metal3 s 0 26604 800 26844 6 la1_data_out[0]
port 148 nsew signal output
rlabel metal3 s 0 34764 800 35004 6 la1_data_out[10]
port 149 nsew signal output
rlabel metal3 s 0 35580 800 35820 6 la1_data_out[11]
port 150 nsew signal output
rlabel metal3 s 0 36396 800 36636 6 la1_data_out[12]
port 151 nsew signal output
rlabel metal3 s 0 37212 800 37452 6 la1_data_out[13]
port 152 nsew signal output
rlabel metal3 s 0 38028 800 38268 6 la1_data_out[14]
port 153 nsew signal output
rlabel metal3 s 0 38844 800 39084 6 la1_data_out[15]
port 154 nsew signal output
rlabel metal3 s 0 39660 800 39900 6 la1_data_out[16]
port 155 nsew signal output
rlabel metal3 s 0 40612 800 40852 6 la1_data_out[17]
port 156 nsew signal output
rlabel metal3 s 0 41428 800 41668 6 la1_data_out[18]
port 157 nsew signal output
rlabel metal3 s 0 42244 800 42484 6 la1_data_out[19]
port 158 nsew signal output
rlabel metal3 s 0 27420 800 27660 6 la1_data_out[1]
port 159 nsew signal output
rlabel metal3 s 0 43060 800 43300 6 la1_data_out[20]
port 160 nsew signal output
rlabel metal3 s 0 43876 800 44116 6 la1_data_out[21]
port 161 nsew signal output
rlabel metal3 s 0 44692 800 44932 6 la1_data_out[22]
port 162 nsew signal output
rlabel metal3 s 0 45508 800 45748 6 la1_data_out[23]
port 163 nsew signal output
rlabel metal3 s 0 46324 800 46564 6 la1_data_out[24]
port 164 nsew signal output
rlabel metal3 s 0 47140 800 47380 6 la1_data_out[25]
port 165 nsew signal output
rlabel metal3 s 0 47956 800 48196 6 la1_data_out[26]
port 166 nsew signal output
rlabel metal3 s 0 48772 800 49012 6 la1_data_out[27]
port 167 nsew signal output
rlabel metal3 s 0 49588 800 49828 6 la1_data_out[28]
port 168 nsew signal output
rlabel metal3 s 0 50404 800 50644 6 la1_data_out[29]
port 169 nsew signal output
rlabel metal3 s 0 28236 800 28476 6 la1_data_out[2]
port 170 nsew signal output
rlabel metal3 s 0 51220 800 51460 6 la1_data_out[30]
port 171 nsew signal output
rlabel metal3 s 0 52036 800 52276 6 la1_data_out[31]
port 172 nsew signal output
rlabel metal3 s 0 29052 800 29292 6 la1_data_out[3]
port 173 nsew signal output
rlabel metal3 s 0 29868 800 30108 6 la1_data_out[4]
port 174 nsew signal output
rlabel metal3 s 0 30684 800 30924 6 la1_data_out[5]
port 175 nsew signal output
rlabel metal3 s 0 31500 800 31740 6 la1_data_out[6]
port 176 nsew signal output
rlabel metal3 s 0 32316 800 32556 6 la1_data_out[7]
port 177 nsew signal output
rlabel metal3 s 0 33132 800 33372 6 la1_data_out[8]
port 178 nsew signal output
rlabel metal3 s 0 33948 800 34188 6 la1_data_out[9]
port 179 nsew signal output
rlabel metal3 s 59200 220 60000 460 6 la1_oenb[0]
port 180 nsew signal input
rlabel metal3 s 59200 7564 60000 7804 6 la1_oenb[10]
port 181 nsew signal input
rlabel metal3 s 59200 8244 60000 8484 6 la1_oenb[11]
port 182 nsew signal input
rlabel metal3 s 59200 9060 60000 9300 6 la1_oenb[12]
port 183 nsew signal input
rlabel metal3 s 59200 9740 60000 9980 6 la1_oenb[13]
port 184 nsew signal input
rlabel metal3 s 59200 10556 60000 10796 6 la1_oenb[14]
port 185 nsew signal input
rlabel metal3 s 59200 11236 60000 11476 6 la1_oenb[15]
port 186 nsew signal input
rlabel metal3 s 59200 12052 60000 12292 6 la1_oenb[16]
port 187 nsew signal input
rlabel metal3 s 59200 12732 60000 12972 6 la1_oenb[17]
port 188 nsew signal input
rlabel metal3 s 59200 13548 60000 13788 6 la1_oenb[18]
port 189 nsew signal input
rlabel metal3 s 59200 14228 60000 14468 6 la1_oenb[19]
port 190 nsew signal input
rlabel metal3 s 59200 900 60000 1140 6 la1_oenb[1]
port 191 nsew signal input
rlabel metal3 s 59200 14908 60000 15148 6 la1_oenb[20]
port 192 nsew signal input
rlabel metal3 s 59200 15724 60000 15964 6 la1_oenb[21]
port 193 nsew signal input
rlabel metal3 s 59200 16404 60000 16644 6 la1_oenb[22]
port 194 nsew signal input
rlabel metal3 s 59200 17220 60000 17460 6 la1_oenb[23]
port 195 nsew signal input
rlabel metal3 s 59200 17900 60000 18140 6 la1_oenb[24]
port 196 nsew signal input
rlabel metal3 s 59200 18716 60000 18956 6 la1_oenb[25]
port 197 nsew signal input
rlabel metal3 s 59200 19396 60000 19636 6 la1_oenb[26]
port 198 nsew signal input
rlabel metal3 s 59200 20212 60000 20452 6 la1_oenb[27]
port 199 nsew signal input
rlabel metal3 s 59200 20892 60000 21132 6 la1_oenb[28]
port 200 nsew signal input
rlabel metal3 s 59200 21572 60000 21812 6 la1_oenb[29]
port 201 nsew signal input
rlabel metal3 s 59200 1580 60000 1820 6 la1_oenb[2]
port 202 nsew signal input
rlabel metal3 s 59200 22388 60000 22628 6 la1_oenb[30]
port 203 nsew signal input
rlabel metal3 s 59200 23068 60000 23308 6 la1_oenb[31]
port 204 nsew signal input
rlabel metal3 s 59200 2396 60000 2636 6 la1_oenb[3]
port 205 nsew signal input
rlabel metal3 s 59200 3076 60000 3316 6 la1_oenb[4]
port 206 nsew signal input
rlabel metal3 s 59200 3892 60000 4132 6 la1_oenb[5]
port 207 nsew signal input
rlabel metal3 s 59200 4572 60000 4812 6 la1_oenb[6]
port 208 nsew signal input
rlabel metal3 s 59200 5388 60000 5628 6 la1_oenb[7]
port 209 nsew signal input
rlabel metal3 s 59200 6068 60000 6308 6 la1_oenb[8]
port 210 nsew signal input
rlabel metal3 s 59200 6884 60000 7124 6 la1_oenb[9]
port 211 nsew signal input
rlabel metal4 s 4208 496 4528 57712 6 vccd1
port 212 nsew power input
rlabel metal4 s 34928 496 35248 57712 6 vccd1
port 212 nsew power input
rlabel metal4 s 19568 496 19888 57712 6 vssd1
port 213 nsew ground input
rlabel metal4 s 50288 496 50608 57712 6 vssd1
port 213 nsew ground input
rlabel metal2 s 1738 59200 1850 60000 6 wb_clk_i
port 214 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 60000 60000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 12332516
string GDS_FILE /openlane/designs/wrapped-vgademo-on-fpga/runs/RUN_2022.03.20_07.24.20/results/finishing/wrapped_vgademo_on_fpga.magic.gds
string GDS_START 1105746
<< end >>

