magic
tech sky130A
magscale 1 2
timestamp 1647850625
<< obsli1 >>
rect 1104 527 58880 57681
<< obsm1 >>
rect 566 416 59418 57860
<< metal2 >>
rect 542 59200 654 60000
rect 1646 59200 1758 60000
rect 2842 59200 2954 60000
rect 3946 59200 4058 60000
rect 5142 59200 5254 60000
rect 6246 59200 6358 60000
rect 7442 59200 7554 60000
rect 8546 59200 8658 60000
rect 9742 59200 9854 60000
rect 10846 59200 10958 60000
rect 12042 59200 12154 60000
rect 13146 59200 13258 60000
rect 14342 59200 14454 60000
rect 15538 59200 15650 60000
rect 16642 59200 16754 60000
rect 17838 59200 17950 60000
rect 18942 59200 19054 60000
rect 20138 59200 20250 60000
rect 21242 59200 21354 60000
rect 22438 59200 22550 60000
rect 23542 59200 23654 60000
rect 24738 59200 24850 60000
rect 25842 59200 25954 60000
rect 27038 59200 27150 60000
rect 28142 59200 28254 60000
rect 29338 59200 29450 60000
rect 30534 59200 30646 60000
rect 31638 59200 31750 60000
rect 32834 59200 32946 60000
rect 33938 59200 34050 60000
rect 35134 59200 35246 60000
rect 36238 59200 36350 60000
rect 37434 59200 37546 60000
rect 38538 59200 38650 60000
rect 39734 59200 39846 60000
rect 40838 59200 40950 60000
rect 42034 59200 42146 60000
rect 43138 59200 43250 60000
rect 44334 59200 44446 60000
rect 45530 59200 45642 60000
rect 46634 59200 46746 60000
rect 47830 59200 47942 60000
rect 48934 59200 49046 60000
rect 50130 59200 50242 60000
rect 51234 59200 51346 60000
rect 52430 59200 52542 60000
rect 53534 59200 53646 60000
rect 54730 59200 54842 60000
rect 55834 59200 55946 60000
rect 57030 59200 57142 60000
rect 58134 59200 58246 60000
rect 59330 59200 59442 60000
rect 4222 0 4334 800
rect 12778 0 12890 800
rect 21334 0 21446 800
rect 29890 0 30002 800
rect 38446 0 38558 800
rect 47002 0 47114 800
rect 55558 0 55670 800
<< obsm2 >>
rect 710 59144 1590 59537
rect 1814 59144 2786 59537
rect 3010 59144 3890 59537
rect 4114 59144 5086 59537
rect 5310 59144 6190 59537
rect 6414 59144 7386 59537
rect 7610 59144 8490 59537
rect 8714 59144 9686 59537
rect 9910 59144 10790 59537
rect 11014 59144 11986 59537
rect 12210 59144 13090 59537
rect 13314 59144 14286 59537
rect 14510 59144 15482 59537
rect 15706 59144 16586 59537
rect 16810 59144 17782 59537
rect 18006 59144 18886 59537
rect 19110 59144 20082 59537
rect 20306 59144 21186 59537
rect 21410 59144 22382 59537
rect 22606 59144 23486 59537
rect 23710 59144 24682 59537
rect 24906 59144 25786 59537
rect 26010 59144 26982 59537
rect 27206 59144 28086 59537
rect 28310 59144 29282 59537
rect 29506 59144 30478 59537
rect 30702 59144 31582 59537
rect 31806 59144 32778 59537
rect 33002 59144 33882 59537
rect 34106 59144 35078 59537
rect 35302 59144 36182 59537
rect 36406 59144 37378 59537
rect 37602 59144 38482 59537
rect 38706 59144 39678 59537
rect 39902 59144 40782 59537
rect 41006 59144 41978 59537
rect 42202 59144 43082 59537
rect 43306 59144 44278 59537
rect 44502 59144 45474 59537
rect 45698 59144 46578 59537
rect 46802 59144 47774 59537
rect 47998 59144 48878 59537
rect 49102 59144 50074 59537
rect 50298 59144 51178 59537
rect 51402 59144 52374 59537
rect 52598 59144 53478 59537
rect 53702 59144 54674 59537
rect 54898 59144 55778 59537
rect 56002 59144 56974 59537
rect 57198 59144 58078 59537
rect 58302 59144 59274 59537
rect 572 856 59412 59144
rect 572 410 4166 856
rect 4390 410 12722 856
rect 12946 410 21278 856
rect 21502 410 29834 856
rect 30058 410 38390 856
rect 38614 410 46946 856
rect 47170 410 55502 856
rect 55726 410 59412 856
<< metal3 >>
rect 0 59380 800 59620
rect 59200 59380 60000 59620
rect 0 58564 800 58804
rect 59200 58700 60000 58940
rect 59200 58020 60000 58260
rect 0 57612 800 57852
rect 59200 57340 60000 57580
rect 0 56796 800 57036
rect 59200 56524 60000 56764
rect 0 55980 800 56220
rect 59200 55844 60000 56084
rect 0 55028 800 55268
rect 59200 55164 60000 55404
rect 0 54212 800 54452
rect 59200 54484 60000 54724
rect 59200 53668 60000 53908
rect 0 53260 800 53500
rect 59200 52988 60000 53228
rect 0 52444 800 52684
rect 59200 52308 60000 52548
rect 0 51628 800 51868
rect 59200 51628 60000 51868
rect 0 50676 800 50916
rect 59200 50812 60000 51052
rect 0 49860 800 50100
rect 59200 50132 60000 50372
rect 59200 49452 60000 49692
rect 0 48908 800 49148
rect 59200 48772 60000 49012
rect 0 48092 800 48332
rect 59200 47956 60000 48196
rect 0 47276 800 47516
rect 59200 47276 60000 47516
rect 0 46324 800 46564
rect 59200 46596 60000 46836
rect 59200 45916 60000 46156
rect 0 45508 800 45748
rect 59200 45100 60000 45340
rect 0 44556 800 44796
rect 59200 44420 60000 44660
rect 0 43740 800 43980
rect 59200 43740 60000 43980
rect 0 42924 800 43164
rect 59200 43060 60000 43300
rect 0 41972 800 42212
rect 59200 42244 60000 42484
rect 59200 41564 60000 41804
rect 0 41156 800 41396
rect 59200 40884 60000 41124
rect 0 40340 800 40580
rect 59200 40204 60000 40444
rect 0 39388 800 39628
rect 59200 39388 60000 39628
rect 0 38572 800 38812
rect 59200 38708 60000 38948
rect 59200 38028 60000 38268
rect 0 37620 800 37860
rect 59200 37348 60000 37588
rect 0 36804 800 37044
rect 59200 36532 60000 36772
rect 0 35988 800 36228
rect 59200 35852 60000 36092
rect 0 35036 800 35276
rect 59200 35172 60000 35412
rect 0 34220 800 34460
rect 59200 34492 60000 34732
rect 59200 33676 60000 33916
rect 0 33268 800 33508
rect 59200 32996 60000 33236
rect 0 32452 800 32692
rect 59200 32316 60000 32556
rect 0 31636 800 31876
rect 59200 31636 60000 31876
rect 0 30684 800 30924
rect 59200 30820 60000 31060
rect 0 29868 800 30108
rect 59200 30140 60000 30380
rect 59200 29460 60000 29700
rect 0 28916 800 29156
rect 59200 28780 60000 29020
rect 0 28100 800 28340
rect 59200 27964 60000 28204
rect 0 27284 800 27524
rect 59200 27284 60000 27524
rect 0 26332 800 26572
rect 59200 26604 60000 26844
rect 59200 25924 60000 26164
rect 0 25516 800 25756
rect 59200 25108 60000 25348
rect 0 24564 800 24804
rect 59200 24428 60000 24668
rect 0 23748 800 23988
rect 59200 23748 60000 23988
rect 0 22932 800 23172
rect 59200 23068 60000 23308
rect 0 21980 800 22220
rect 59200 22252 60000 22492
rect 59200 21572 60000 21812
rect 0 21164 800 21404
rect 59200 20892 60000 21132
rect 0 20348 800 20588
rect 59200 20212 60000 20452
rect 0 19396 800 19636
rect 59200 19396 60000 19636
rect 0 18580 800 18820
rect 59200 18716 60000 18956
rect 59200 18036 60000 18276
rect 0 17628 800 17868
rect 59200 17356 60000 17596
rect 0 16812 800 17052
rect 59200 16540 60000 16780
rect 0 15996 800 16236
rect 59200 15860 60000 16100
rect 0 15044 800 15284
rect 59200 15180 60000 15420
rect 0 14228 800 14468
rect 59200 14500 60000 14740
rect 59200 13684 60000 13924
rect 0 13276 800 13516
rect 59200 13004 60000 13244
rect 0 12460 800 12700
rect 59200 12324 60000 12564
rect 0 11644 800 11884
rect 59200 11644 60000 11884
rect 0 10692 800 10932
rect 59200 10828 60000 11068
rect 0 9876 800 10116
rect 59200 10148 60000 10388
rect 59200 9468 60000 9708
rect 0 8924 800 9164
rect 59200 8788 60000 9028
rect 0 8108 800 8348
rect 59200 7972 60000 8212
rect 0 7292 800 7532
rect 59200 7292 60000 7532
rect 0 6340 800 6580
rect 59200 6612 60000 6852
rect 59200 5932 60000 6172
rect 0 5524 800 5764
rect 59200 5116 60000 5356
rect 0 4572 800 4812
rect 59200 4436 60000 4676
rect 0 3756 800 3996
rect 59200 3756 60000 3996
rect 0 2940 800 3180
rect 59200 3076 60000 3316
rect 0 1988 800 2228
rect 59200 2260 60000 2500
rect 59200 1580 60000 1820
rect 0 1172 800 1412
rect 59200 900 60000 1140
rect 0 356 800 596
rect 59200 220 60000 460
<< obsm3 >>
rect 880 59300 59120 59533
rect 800 59020 59200 59300
rect 800 58884 59120 59020
rect 880 58620 59120 58884
rect 880 58484 59200 58620
rect 800 58340 59200 58484
rect 800 57940 59120 58340
rect 800 57932 59200 57940
rect 880 57660 59200 57932
rect 880 57532 59120 57660
rect 800 57260 59120 57532
rect 800 57116 59200 57260
rect 880 56844 59200 57116
rect 880 56716 59120 56844
rect 800 56444 59120 56716
rect 800 56300 59200 56444
rect 880 56164 59200 56300
rect 880 55900 59120 56164
rect 800 55764 59120 55900
rect 800 55484 59200 55764
rect 800 55348 59120 55484
rect 880 55084 59120 55348
rect 880 54948 59200 55084
rect 800 54804 59200 54948
rect 800 54532 59120 54804
rect 880 54404 59120 54532
rect 880 54132 59200 54404
rect 800 53988 59200 54132
rect 800 53588 59120 53988
rect 800 53580 59200 53588
rect 880 53308 59200 53580
rect 880 53180 59120 53308
rect 800 52908 59120 53180
rect 800 52764 59200 52908
rect 880 52628 59200 52764
rect 880 52364 59120 52628
rect 800 52228 59120 52364
rect 800 51948 59200 52228
rect 880 51548 59120 51948
rect 800 51132 59200 51548
rect 800 50996 59120 51132
rect 880 50732 59120 50996
rect 880 50596 59200 50732
rect 800 50452 59200 50596
rect 800 50180 59120 50452
rect 880 50052 59120 50180
rect 880 49780 59200 50052
rect 800 49772 59200 49780
rect 800 49372 59120 49772
rect 800 49228 59200 49372
rect 880 49092 59200 49228
rect 880 48828 59120 49092
rect 800 48692 59120 48828
rect 800 48412 59200 48692
rect 880 48276 59200 48412
rect 880 48012 59120 48276
rect 800 47876 59120 48012
rect 800 47596 59200 47876
rect 880 47196 59120 47596
rect 800 46916 59200 47196
rect 800 46644 59120 46916
rect 880 46516 59120 46644
rect 880 46244 59200 46516
rect 800 46236 59200 46244
rect 800 45836 59120 46236
rect 800 45828 59200 45836
rect 880 45428 59200 45828
rect 800 45420 59200 45428
rect 800 45020 59120 45420
rect 800 44876 59200 45020
rect 880 44740 59200 44876
rect 880 44476 59120 44740
rect 800 44340 59120 44476
rect 800 44060 59200 44340
rect 880 43660 59120 44060
rect 800 43380 59200 43660
rect 800 43244 59120 43380
rect 880 42980 59120 43244
rect 880 42844 59200 42980
rect 800 42564 59200 42844
rect 800 42292 59120 42564
rect 880 42164 59120 42292
rect 880 41892 59200 42164
rect 800 41884 59200 41892
rect 800 41484 59120 41884
rect 800 41476 59200 41484
rect 880 41204 59200 41476
rect 880 41076 59120 41204
rect 800 40804 59120 41076
rect 800 40660 59200 40804
rect 880 40524 59200 40660
rect 880 40260 59120 40524
rect 800 40124 59120 40260
rect 800 39708 59200 40124
rect 880 39308 59120 39708
rect 800 39028 59200 39308
rect 800 38892 59120 39028
rect 880 38628 59120 38892
rect 880 38492 59200 38628
rect 800 38348 59200 38492
rect 800 37948 59120 38348
rect 800 37940 59200 37948
rect 880 37668 59200 37940
rect 880 37540 59120 37668
rect 800 37268 59120 37540
rect 800 37124 59200 37268
rect 880 36852 59200 37124
rect 880 36724 59120 36852
rect 800 36452 59120 36724
rect 800 36308 59200 36452
rect 880 36172 59200 36308
rect 880 35908 59120 36172
rect 800 35772 59120 35908
rect 800 35492 59200 35772
rect 800 35356 59120 35492
rect 880 35092 59120 35356
rect 880 34956 59200 35092
rect 800 34812 59200 34956
rect 800 34540 59120 34812
rect 880 34412 59120 34540
rect 880 34140 59200 34412
rect 800 33996 59200 34140
rect 800 33596 59120 33996
rect 800 33588 59200 33596
rect 880 33316 59200 33588
rect 880 33188 59120 33316
rect 800 32916 59120 33188
rect 800 32772 59200 32916
rect 880 32636 59200 32772
rect 880 32372 59120 32636
rect 800 32236 59120 32372
rect 800 31956 59200 32236
rect 880 31556 59120 31956
rect 800 31140 59200 31556
rect 800 31004 59120 31140
rect 880 30740 59120 31004
rect 880 30604 59200 30740
rect 800 30460 59200 30604
rect 800 30188 59120 30460
rect 880 30060 59120 30188
rect 880 29788 59200 30060
rect 800 29780 59200 29788
rect 800 29380 59120 29780
rect 800 29236 59200 29380
rect 880 29100 59200 29236
rect 880 28836 59120 29100
rect 800 28700 59120 28836
rect 800 28420 59200 28700
rect 880 28284 59200 28420
rect 880 28020 59120 28284
rect 800 27884 59120 28020
rect 800 27604 59200 27884
rect 880 27204 59120 27604
rect 800 26924 59200 27204
rect 800 26652 59120 26924
rect 880 26524 59120 26652
rect 880 26252 59200 26524
rect 800 26244 59200 26252
rect 800 25844 59120 26244
rect 800 25836 59200 25844
rect 880 25436 59200 25836
rect 800 25428 59200 25436
rect 800 25028 59120 25428
rect 800 24884 59200 25028
rect 880 24748 59200 24884
rect 880 24484 59120 24748
rect 800 24348 59120 24484
rect 800 24068 59200 24348
rect 880 23668 59120 24068
rect 800 23388 59200 23668
rect 800 23252 59120 23388
rect 880 22988 59120 23252
rect 880 22852 59200 22988
rect 800 22572 59200 22852
rect 800 22300 59120 22572
rect 880 22172 59120 22300
rect 880 21900 59200 22172
rect 800 21892 59200 21900
rect 800 21492 59120 21892
rect 800 21484 59200 21492
rect 880 21212 59200 21484
rect 880 21084 59120 21212
rect 800 20812 59120 21084
rect 800 20668 59200 20812
rect 880 20532 59200 20668
rect 880 20268 59120 20532
rect 800 20132 59120 20268
rect 800 19716 59200 20132
rect 880 19316 59120 19716
rect 800 19036 59200 19316
rect 800 18900 59120 19036
rect 880 18636 59120 18900
rect 880 18500 59200 18636
rect 800 18356 59200 18500
rect 800 17956 59120 18356
rect 800 17948 59200 17956
rect 880 17676 59200 17948
rect 880 17548 59120 17676
rect 800 17276 59120 17548
rect 800 17132 59200 17276
rect 880 16860 59200 17132
rect 880 16732 59120 16860
rect 800 16460 59120 16732
rect 800 16316 59200 16460
rect 880 16180 59200 16316
rect 880 15916 59120 16180
rect 800 15780 59120 15916
rect 800 15500 59200 15780
rect 800 15364 59120 15500
rect 880 15100 59120 15364
rect 880 14964 59200 15100
rect 800 14820 59200 14964
rect 800 14548 59120 14820
rect 880 14420 59120 14548
rect 880 14148 59200 14420
rect 800 14004 59200 14148
rect 800 13604 59120 14004
rect 800 13596 59200 13604
rect 880 13324 59200 13596
rect 880 13196 59120 13324
rect 800 12924 59120 13196
rect 800 12780 59200 12924
rect 880 12644 59200 12780
rect 880 12380 59120 12644
rect 800 12244 59120 12380
rect 800 11964 59200 12244
rect 880 11564 59120 11964
rect 800 11148 59200 11564
rect 800 11012 59120 11148
rect 880 10748 59120 11012
rect 880 10612 59200 10748
rect 800 10468 59200 10612
rect 800 10196 59120 10468
rect 880 10068 59120 10196
rect 880 9796 59200 10068
rect 800 9788 59200 9796
rect 800 9388 59120 9788
rect 800 9244 59200 9388
rect 880 9108 59200 9244
rect 880 8844 59120 9108
rect 800 8708 59120 8844
rect 800 8428 59200 8708
rect 880 8292 59200 8428
rect 880 8028 59120 8292
rect 800 7892 59120 8028
rect 800 7612 59200 7892
rect 880 7212 59120 7612
rect 800 6932 59200 7212
rect 800 6660 59120 6932
rect 880 6532 59120 6660
rect 880 6260 59200 6532
rect 800 6252 59200 6260
rect 800 5852 59120 6252
rect 800 5844 59200 5852
rect 880 5444 59200 5844
rect 800 5436 59200 5444
rect 800 5036 59120 5436
rect 800 4892 59200 5036
rect 880 4756 59200 4892
rect 880 4492 59120 4756
rect 800 4356 59120 4492
rect 800 4076 59200 4356
rect 880 3676 59120 4076
rect 800 3396 59200 3676
rect 800 3260 59120 3396
rect 880 2996 59120 3260
rect 880 2860 59200 2996
rect 800 2580 59200 2860
rect 800 2308 59120 2580
rect 880 2180 59120 2308
rect 880 1908 59200 2180
rect 800 1900 59200 1908
rect 800 1500 59120 1900
rect 800 1492 59200 1500
rect 880 1220 59200 1492
rect 880 1092 59120 1220
rect 800 820 59120 1092
rect 800 676 59200 820
rect 880 540 59200 676
rect 880 511 59120 540
<< metal4 >>
rect 4208 496 4528 57712
rect 19568 496 19888 57712
rect 34928 496 35248 57712
rect 50288 496 50608 57712
<< obsm4 >>
rect 3923 3979 4128 56677
rect 4608 3979 19488 56677
rect 19968 3979 34848 56677
rect 35328 3979 36741 56677
<< labels >>
rlabel metal2 s 542 59200 654 60000 6 active
port 1 nsew signal input
rlabel metal2 s 2842 59200 2954 60000 6 io_in[0]
port 2 nsew signal input
rlabel metal2 s 14342 59200 14454 60000 6 io_in[10]
port 3 nsew signal input
rlabel metal2 s 15538 59200 15650 60000 6 io_in[11]
port 4 nsew signal input
rlabel metal2 s 16642 59200 16754 60000 6 io_in[12]
port 5 nsew signal input
rlabel metal2 s 17838 59200 17950 60000 6 io_in[13]
port 6 nsew signal input
rlabel metal2 s 18942 59200 19054 60000 6 io_in[14]
port 7 nsew signal input
rlabel metal2 s 20138 59200 20250 60000 6 io_in[15]
port 8 nsew signal input
rlabel metal2 s 21242 59200 21354 60000 6 io_in[16]
port 9 nsew signal input
rlabel metal2 s 22438 59200 22550 60000 6 io_in[17]
port 10 nsew signal input
rlabel metal2 s 23542 59200 23654 60000 6 io_in[18]
port 11 nsew signal input
rlabel metal2 s 24738 59200 24850 60000 6 io_in[19]
port 12 nsew signal input
rlabel metal2 s 3946 59200 4058 60000 6 io_in[1]
port 13 nsew signal input
rlabel metal2 s 25842 59200 25954 60000 6 io_in[20]
port 14 nsew signal input
rlabel metal2 s 27038 59200 27150 60000 6 io_in[21]
port 15 nsew signal input
rlabel metal2 s 28142 59200 28254 60000 6 io_in[22]
port 16 nsew signal input
rlabel metal2 s 29338 59200 29450 60000 6 io_in[23]
port 17 nsew signal input
rlabel metal2 s 30534 59200 30646 60000 6 io_in[24]
port 18 nsew signal input
rlabel metal2 s 31638 59200 31750 60000 6 io_in[25]
port 19 nsew signal input
rlabel metal2 s 32834 59200 32946 60000 6 io_in[26]
port 20 nsew signal input
rlabel metal2 s 33938 59200 34050 60000 6 io_in[27]
port 21 nsew signal input
rlabel metal2 s 35134 59200 35246 60000 6 io_in[28]
port 22 nsew signal input
rlabel metal2 s 36238 59200 36350 60000 6 io_in[29]
port 23 nsew signal input
rlabel metal2 s 5142 59200 5254 60000 6 io_in[2]
port 24 nsew signal input
rlabel metal2 s 37434 59200 37546 60000 6 io_in[30]
port 25 nsew signal input
rlabel metal2 s 38538 59200 38650 60000 6 io_in[31]
port 26 nsew signal input
rlabel metal2 s 39734 59200 39846 60000 6 io_in[32]
port 27 nsew signal input
rlabel metal2 s 40838 59200 40950 60000 6 io_in[33]
port 28 nsew signal input
rlabel metal2 s 42034 59200 42146 60000 6 io_in[34]
port 29 nsew signal input
rlabel metal2 s 43138 59200 43250 60000 6 io_in[35]
port 30 nsew signal input
rlabel metal2 s 44334 59200 44446 60000 6 io_in[36]
port 31 nsew signal input
rlabel metal2 s 45530 59200 45642 60000 6 io_in[37]
port 32 nsew signal input
rlabel metal2 s 6246 59200 6358 60000 6 io_in[3]
port 33 nsew signal input
rlabel metal2 s 7442 59200 7554 60000 6 io_in[4]
port 34 nsew signal input
rlabel metal2 s 8546 59200 8658 60000 6 io_in[5]
port 35 nsew signal input
rlabel metal2 s 9742 59200 9854 60000 6 io_in[6]
port 36 nsew signal input
rlabel metal2 s 10846 59200 10958 60000 6 io_in[7]
port 37 nsew signal input
rlabel metal2 s 12042 59200 12154 60000 6 io_in[8]
port 38 nsew signal input
rlabel metal2 s 13146 59200 13258 60000 6 io_in[9]
port 39 nsew signal input
rlabel metal3 s 59200 23068 60000 23308 6 io_oeb[0]
port 40 nsew signal output
rlabel metal3 s 59200 30140 60000 30380 6 io_oeb[10]
port 41 nsew signal output
rlabel metal3 s 59200 30820 60000 31060 6 io_oeb[11]
port 42 nsew signal output
rlabel metal3 s 59200 31636 60000 31876 6 io_oeb[12]
port 43 nsew signal output
rlabel metal3 s 59200 32316 60000 32556 6 io_oeb[13]
port 44 nsew signal output
rlabel metal3 s 59200 32996 60000 33236 6 io_oeb[14]
port 45 nsew signal output
rlabel metal3 s 59200 33676 60000 33916 6 io_oeb[15]
port 46 nsew signal output
rlabel metal3 s 59200 34492 60000 34732 6 io_oeb[16]
port 47 nsew signal output
rlabel metal3 s 59200 35172 60000 35412 6 io_oeb[17]
port 48 nsew signal output
rlabel metal3 s 59200 35852 60000 36092 6 io_oeb[18]
port 49 nsew signal output
rlabel metal3 s 59200 36532 60000 36772 6 io_oeb[19]
port 50 nsew signal output
rlabel metal3 s 59200 23748 60000 23988 6 io_oeb[1]
port 51 nsew signal output
rlabel metal3 s 59200 37348 60000 37588 6 io_oeb[20]
port 52 nsew signal output
rlabel metal3 s 59200 38028 60000 38268 6 io_oeb[21]
port 53 nsew signal output
rlabel metal3 s 59200 38708 60000 38948 6 io_oeb[22]
port 54 nsew signal output
rlabel metal3 s 59200 39388 60000 39628 6 io_oeb[23]
port 55 nsew signal output
rlabel metal3 s 59200 40204 60000 40444 6 io_oeb[24]
port 56 nsew signal output
rlabel metal3 s 59200 40884 60000 41124 6 io_oeb[25]
port 57 nsew signal output
rlabel metal3 s 59200 41564 60000 41804 6 io_oeb[26]
port 58 nsew signal output
rlabel metal3 s 59200 42244 60000 42484 6 io_oeb[27]
port 59 nsew signal output
rlabel metal3 s 59200 43060 60000 43300 6 io_oeb[28]
port 60 nsew signal output
rlabel metal3 s 59200 43740 60000 43980 6 io_oeb[29]
port 61 nsew signal output
rlabel metal3 s 59200 24428 60000 24668 6 io_oeb[2]
port 62 nsew signal output
rlabel metal3 s 59200 44420 60000 44660 6 io_oeb[30]
port 63 nsew signal output
rlabel metal3 s 59200 45100 60000 45340 6 io_oeb[31]
port 64 nsew signal output
rlabel metal3 s 59200 45916 60000 46156 6 io_oeb[32]
port 65 nsew signal output
rlabel metal3 s 59200 46596 60000 46836 6 io_oeb[33]
port 66 nsew signal output
rlabel metal3 s 59200 47276 60000 47516 6 io_oeb[34]
port 67 nsew signal output
rlabel metal3 s 59200 47956 60000 48196 6 io_oeb[35]
port 68 nsew signal output
rlabel metal3 s 59200 48772 60000 49012 6 io_oeb[36]
port 69 nsew signal output
rlabel metal3 s 59200 49452 60000 49692 6 io_oeb[37]
port 70 nsew signal output
rlabel metal3 s 59200 25108 60000 25348 6 io_oeb[3]
port 71 nsew signal output
rlabel metal3 s 59200 25924 60000 26164 6 io_oeb[4]
port 72 nsew signal output
rlabel metal3 s 59200 26604 60000 26844 6 io_oeb[5]
port 73 nsew signal output
rlabel metal3 s 59200 27284 60000 27524 6 io_oeb[6]
port 74 nsew signal output
rlabel metal3 s 59200 27964 60000 28204 6 io_oeb[7]
port 75 nsew signal output
rlabel metal3 s 59200 28780 60000 29020 6 io_oeb[8]
port 76 nsew signal output
rlabel metal3 s 59200 29460 60000 29700 6 io_oeb[9]
port 77 nsew signal output
rlabel metal3 s 59200 50132 60000 50372 6 io_out[0]
port 78 nsew signal output
rlabel metal3 s 59200 53668 60000 53908 6 io_out[10]
port 79 nsew signal output
rlabel metal3 s 0 55980 800 56220 6 io_out[11]
port 80 nsew signal output
rlabel metal3 s 59200 54484 60000 54724 6 io_out[12]
port 81 nsew signal output
rlabel metal2 s 51234 59200 51346 60000 6 io_out[13]
port 82 nsew signal output
rlabel metal3 s 0 56796 800 57036 6 io_out[14]
port 83 nsew signal output
rlabel metal2 s 52430 59200 52542 60000 6 io_out[15]
port 84 nsew signal output
rlabel metal2 s 12778 0 12890 800 6 io_out[16]
port 85 nsew signal output
rlabel metal3 s 59200 55164 60000 55404 6 io_out[17]
port 86 nsew signal output
rlabel metal3 s 59200 55844 60000 56084 6 io_out[18]
port 87 nsew signal output
rlabel metal2 s 21334 0 21446 800 6 io_out[19]
port 88 nsew signal output
rlabel metal3 s 59200 50812 60000 51052 6 io_out[1]
port 89 nsew signal output
rlabel metal3 s 59200 56524 60000 56764 6 io_out[20]
port 90 nsew signal output
rlabel metal2 s 53534 59200 53646 60000 6 io_out[21]
port 91 nsew signal output
rlabel metal3 s 59200 57340 60000 57580 6 io_out[22]
port 92 nsew signal output
rlabel metal2 s 29890 0 30002 800 6 io_out[23]
port 93 nsew signal output
rlabel metal2 s 54730 59200 54842 60000 6 io_out[24]
port 94 nsew signal output
rlabel metal3 s 0 57612 800 57852 6 io_out[25]
port 95 nsew signal output
rlabel metal2 s 55834 59200 55946 60000 6 io_out[26]
port 96 nsew signal output
rlabel metal3 s 0 58564 800 58804 6 io_out[27]
port 97 nsew signal output
rlabel metal2 s 57030 59200 57142 60000 6 io_out[28]
port 98 nsew signal output
rlabel metal3 s 59200 58020 60000 58260 6 io_out[29]
port 99 nsew signal output
rlabel metal2 s 46634 59200 46746 60000 6 io_out[2]
port 100 nsew signal output
rlabel metal2 s 58134 59200 58246 60000 6 io_out[30]
port 101 nsew signal output
rlabel metal3 s 59200 58700 60000 58940 6 io_out[31]
port 102 nsew signal output
rlabel metal2 s 38446 0 38558 800 6 io_out[32]
port 103 nsew signal output
rlabel metal2 s 47002 0 47114 800 6 io_out[33]
port 104 nsew signal output
rlabel metal2 s 59330 59200 59442 60000 6 io_out[34]
port 105 nsew signal output
rlabel metal3 s 59200 59380 60000 59620 6 io_out[35]
port 106 nsew signal output
rlabel metal3 s 0 59380 800 59620 6 io_out[36]
port 107 nsew signal output
rlabel metal2 s 55558 0 55670 800 6 io_out[37]
port 108 nsew signal output
rlabel metal3 s 59200 51628 60000 51868 6 io_out[3]
port 109 nsew signal output
rlabel metal2 s 47830 59200 47942 60000 6 io_out[4]
port 110 nsew signal output
rlabel metal2 s 48934 59200 49046 60000 6 io_out[5]
port 111 nsew signal output
rlabel metal3 s 59200 52308 60000 52548 6 io_out[6]
port 112 nsew signal output
rlabel metal2 s 4222 0 4334 800 6 io_out[7]
port 113 nsew signal output
rlabel metal2 s 50130 59200 50242 60000 6 io_out[8]
port 114 nsew signal output
rlabel metal3 s 59200 52988 60000 53228 6 io_out[9]
port 115 nsew signal output
rlabel metal3 s 0 356 800 596 6 la1_data_in[0]
port 116 nsew signal input
rlabel metal3 s 0 8924 800 9164 6 la1_data_in[10]
port 117 nsew signal input
rlabel metal3 s 0 9876 800 10116 6 la1_data_in[11]
port 118 nsew signal input
rlabel metal3 s 0 10692 800 10932 6 la1_data_in[12]
port 119 nsew signal input
rlabel metal3 s 0 11644 800 11884 6 la1_data_in[13]
port 120 nsew signal input
rlabel metal3 s 0 12460 800 12700 6 la1_data_in[14]
port 121 nsew signal input
rlabel metal3 s 0 13276 800 13516 6 la1_data_in[15]
port 122 nsew signal input
rlabel metal3 s 0 14228 800 14468 6 la1_data_in[16]
port 123 nsew signal input
rlabel metal3 s 0 15044 800 15284 6 la1_data_in[17]
port 124 nsew signal input
rlabel metal3 s 0 15996 800 16236 6 la1_data_in[18]
port 125 nsew signal input
rlabel metal3 s 0 16812 800 17052 6 la1_data_in[19]
port 126 nsew signal input
rlabel metal3 s 0 1172 800 1412 6 la1_data_in[1]
port 127 nsew signal input
rlabel metal3 s 0 17628 800 17868 6 la1_data_in[20]
port 128 nsew signal input
rlabel metal3 s 0 18580 800 18820 6 la1_data_in[21]
port 129 nsew signal input
rlabel metal3 s 0 19396 800 19636 6 la1_data_in[22]
port 130 nsew signal input
rlabel metal3 s 0 20348 800 20588 6 la1_data_in[23]
port 131 nsew signal input
rlabel metal3 s 0 21164 800 21404 6 la1_data_in[24]
port 132 nsew signal input
rlabel metal3 s 0 21980 800 22220 6 la1_data_in[25]
port 133 nsew signal input
rlabel metal3 s 0 22932 800 23172 6 la1_data_in[26]
port 134 nsew signal input
rlabel metal3 s 0 23748 800 23988 6 la1_data_in[27]
port 135 nsew signal input
rlabel metal3 s 0 24564 800 24804 6 la1_data_in[28]
port 136 nsew signal input
rlabel metal3 s 0 25516 800 25756 6 la1_data_in[29]
port 137 nsew signal input
rlabel metal3 s 0 1988 800 2228 6 la1_data_in[2]
port 138 nsew signal input
rlabel metal3 s 0 26332 800 26572 6 la1_data_in[30]
port 139 nsew signal input
rlabel metal3 s 0 27284 800 27524 6 la1_data_in[31]
port 140 nsew signal input
rlabel metal3 s 0 2940 800 3180 6 la1_data_in[3]
port 141 nsew signal input
rlabel metal3 s 0 3756 800 3996 6 la1_data_in[4]
port 142 nsew signal input
rlabel metal3 s 0 4572 800 4812 6 la1_data_in[5]
port 143 nsew signal input
rlabel metal3 s 0 5524 800 5764 6 la1_data_in[6]
port 144 nsew signal input
rlabel metal3 s 0 6340 800 6580 6 la1_data_in[7]
port 145 nsew signal input
rlabel metal3 s 0 7292 800 7532 6 la1_data_in[8]
port 146 nsew signal input
rlabel metal3 s 0 8108 800 8348 6 la1_data_in[9]
port 147 nsew signal input
rlabel metal3 s 0 28100 800 28340 6 la1_data_out[0]
port 148 nsew signal output
rlabel metal3 s 0 36804 800 37044 6 la1_data_out[10]
port 149 nsew signal output
rlabel metal3 s 0 37620 800 37860 6 la1_data_out[11]
port 150 nsew signal output
rlabel metal3 s 0 38572 800 38812 6 la1_data_out[12]
port 151 nsew signal output
rlabel metal3 s 0 39388 800 39628 6 la1_data_out[13]
port 152 nsew signal output
rlabel metal3 s 0 40340 800 40580 6 la1_data_out[14]
port 153 nsew signal output
rlabel metal3 s 0 41156 800 41396 6 la1_data_out[15]
port 154 nsew signal output
rlabel metal3 s 0 41972 800 42212 6 la1_data_out[16]
port 155 nsew signal output
rlabel metal3 s 0 42924 800 43164 6 la1_data_out[17]
port 156 nsew signal output
rlabel metal3 s 0 43740 800 43980 6 la1_data_out[18]
port 157 nsew signal output
rlabel metal3 s 0 44556 800 44796 6 la1_data_out[19]
port 158 nsew signal output
rlabel metal3 s 0 28916 800 29156 6 la1_data_out[1]
port 159 nsew signal output
rlabel metal3 s 0 45508 800 45748 6 la1_data_out[20]
port 160 nsew signal output
rlabel metal3 s 0 46324 800 46564 6 la1_data_out[21]
port 161 nsew signal output
rlabel metal3 s 0 47276 800 47516 6 la1_data_out[22]
port 162 nsew signal output
rlabel metal3 s 0 48092 800 48332 6 la1_data_out[23]
port 163 nsew signal output
rlabel metal3 s 0 48908 800 49148 6 la1_data_out[24]
port 164 nsew signal output
rlabel metal3 s 0 49860 800 50100 6 la1_data_out[25]
port 165 nsew signal output
rlabel metal3 s 0 50676 800 50916 6 la1_data_out[26]
port 166 nsew signal output
rlabel metal3 s 0 51628 800 51868 6 la1_data_out[27]
port 167 nsew signal output
rlabel metal3 s 0 52444 800 52684 6 la1_data_out[28]
port 168 nsew signal output
rlabel metal3 s 0 53260 800 53500 6 la1_data_out[29]
port 169 nsew signal output
rlabel metal3 s 0 29868 800 30108 6 la1_data_out[2]
port 170 nsew signal output
rlabel metal3 s 0 54212 800 54452 6 la1_data_out[30]
port 171 nsew signal output
rlabel metal3 s 0 55028 800 55268 6 la1_data_out[31]
port 172 nsew signal output
rlabel metal3 s 0 30684 800 30924 6 la1_data_out[3]
port 173 nsew signal output
rlabel metal3 s 0 31636 800 31876 6 la1_data_out[4]
port 174 nsew signal output
rlabel metal3 s 0 32452 800 32692 6 la1_data_out[5]
port 175 nsew signal output
rlabel metal3 s 0 33268 800 33508 6 la1_data_out[6]
port 176 nsew signal output
rlabel metal3 s 0 34220 800 34460 6 la1_data_out[7]
port 177 nsew signal output
rlabel metal3 s 0 35036 800 35276 6 la1_data_out[8]
port 178 nsew signal output
rlabel metal3 s 0 35988 800 36228 6 la1_data_out[9]
port 179 nsew signal output
rlabel metal3 s 59200 220 60000 460 6 la1_oenb[0]
port 180 nsew signal input
rlabel metal3 s 59200 7292 60000 7532 6 la1_oenb[10]
port 181 nsew signal input
rlabel metal3 s 59200 7972 60000 8212 6 la1_oenb[11]
port 182 nsew signal input
rlabel metal3 s 59200 8788 60000 9028 6 la1_oenb[12]
port 183 nsew signal input
rlabel metal3 s 59200 9468 60000 9708 6 la1_oenb[13]
port 184 nsew signal input
rlabel metal3 s 59200 10148 60000 10388 6 la1_oenb[14]
port 185 nsew signal input
rlabel metal3 s 59200 10828 60000 11068 6 la1_oenb[15]
port 186 nsew signal input
rlabel metal3 s 59200 11644 60000 11884 6 la1_oenb[16]
port 187 nsew signal input
rlabel metal3 s 59200 12324 60000 12564 6 la1_oenb[17]
port 188 nsew signal input
rlabel metal3 s 59200 13004 60000 13244 6 la1_oenb[18]
port 189 nsew signal input
rlabel metal3 s 59200 13684 60000 13924 6 la1_oenb[19]
port 190 nsew signal input
rlabel metal3 s 59200 900 60000 1140 6 la1_oenb[1]
port 191 nsew signal input
rlabel metal3 s 59200 14500 60000 14740 6 la1_oenb[20]
port 192 nsew signal input
rlabel metal3 s 59200 15180 60000 15420 6 la1_oenb[21]
port 193 nsew signal input
rlabel metal3 s 59200 15860 60000 16100 6 la1_oenb[22]
port 194 nsew signal input
rlabel metal3 s 59200 16540 60000 16780 6 la1_oenb[23]
port 195 nsew signal input
rlabel metal3 s 59200 17356 60000 17596 6 la1_oenb[24]
port 196 nsew signal input
rlabel metal3 s 59200 18036 60000 18276 6 la1_oenb[25]
port 197 nsew signal input
rlabel metal3 s 59200 18716 60000 18956 6 la1_oenb[26]
port 198 nsew signal input
rlabel metal3 s 59200 19396 60000 19636 6 la1_oenb[27]
port 199 nsew signal input
rlabel metal3 s 59200 20212 60000 20452 6 la1_oenb[28]
port 200 nsew signal input
rlabel metal3 s 59200 20892 60000 21132 6 la1_oenb[29]
port 201 nsew signal input
rlabel metal3 s 59200 1580 60000 1820 6 la1_oenb[2]
port 202 nsew signal input
rlabel metal3 s 59200 21572 60000 21812 6 la1_oenb[30]
port 203 nsew signal input
rlabel metal3 s 59200 22252 60000 22492 6 la1_oenb[31]
port 204 nsew signal input
rlabel metal3 s 59200 2260 60000 2500 6 la1_oenb[3]
port 205 nsew signal input
rlabel metal3 s 59200 3076 60000 3316 6 la1_oenb[4]
port 206 nsew signal input
rlabel metal3 s 59200 3756 60000 3996 6 la1_oenb[5]
port 207 nsew signal input
rlabel metal3 s 59200 4436 60000 4676 6 la1_oenb[6]
port 208 nsew signal input
rlabel metal3 s 59200 5116 60000 5356 6 la1_oenb[7]
port 209 nsew signal input
rlabel metal3 s 59200 5932 60000 6172 6 la1_oenb[8]
port 210 nsew signal input
rlabel metal3 s 59200 6612 60000 6852 6 la1_oenb[9]
port 211 nsew signal input
rlabel metal4 s 4208 496 4528 57712 6 vccd1
port 212 nsew power input
rlabel metal4 s 34928 496 35248 57712 6 vccd1
port 212 nsew power input
rlabel metal4 s 19568 496 19888 57712 6 vssd1
port 213 nsew ground input
rlabel metal4 s 50288 496 50608 57712 6 vssd1
port 213 nsew ground input
rlabel metal2 s 1646 59200 1758 60000 6 wb_clk_i
port 214 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 60000 60000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 12723636
string GDS_FILE /openlane/designs/wrapped-vgademo-on-fpga/runs/RUN_2022.03.21_08.12.07/results/finishing/wrapped_vgademo_on_fpga.magic.gds
string GDS_START 1087710
<< end >>

