VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_vgademo_on_fpga
  CLASS BLOCK ;
  FOREIGN wrapped_vgademo_on_fpga ;
  ORIGIN 0.000 0.000 ;
  SIZE 300.000 BY 300.000 ;
  PIN active
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.710 296.000 3.270 300.000 ;
    END
  END active
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.750 296.000 14.310 300.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.330 296.000 70.890 300.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.850 296.000 76.410 300.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.830 296.000 82.390 300.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.350 296.000 87.910 300.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.870 296.000 93.430 300.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.850 296.000 99.410 300.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.370 296.000 104.930 300.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.890 296.000 110.450 300.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.870 296.000 116.430 300.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.390 296.000 121.950 300.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.270 296.000 19.830 300.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.910 296.000 127.470 300.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.430 296.000 132.990 300.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.410 296.000 138.970 300.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.930 296.000 144.490 300.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.450 296.000 150.010 300.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.430 296.000 155.990 300.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.950 296.000 161.510 300.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.470 296.000 167.030 300.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.450 296.000 173.010 300.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.970 296.000 178.530 300.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.250 296.000 25.810 300.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.490 296.000 184.050 300.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.010 296.000 189.570 300.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.990 296.000 195.550 300.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.510 296.000 201.070 300.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.030 296.000 206.590 300.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.010 296.000 212.570 300.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.530 296.000 218.090 300.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.050 296.000 223.610 300.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.770 296.000 31.330 300.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.290 296.000 36.850 300.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.270 296.000 42.830 300.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.790 296.000 48.350 300.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.310 296.000 53.870 300.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.290 296.000 59.850 300.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.810 296.000 65.370 300.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 122.140 300.000 123.340 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 160.220 300.000 161.420 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 164.300 300.000 165.500 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 167.700 300.000 168.900 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 171.780 300.000 172.980 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 175.180 300.000 176.380 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 179.260 300.000 180.460 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 182.660 300.000 183.860 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 186.740 300.000 187.940 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 190.820 300.000 192.020 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 194.220 300.000 195.420 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 126.220 300.000 127.420 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 198.300 300.000 199.500 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 201.700 300.000 202.900 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 205.780 300.000 206.980 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 209.860 300.000 211.060 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 213.260 300.000 214.460 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 217.340 300.000 218.540 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 220.740 300.000 221.940 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 224.820 300.000 226.020 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 228.220 300.000 229.420 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 232.300 300.000 233.500 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 129.620 300.000 130.820 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 236.380 300.000 237.580 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 239.780 300.000 240.980 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 243.860 300.000 245.060 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 247.260 300.000 248.460 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 251.340 300.000 252.540 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 255.420 300.000 256.620 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 258.820 300.000 260.020 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 262.900 300.000 264.100 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 133.700 300.000 134.900 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 137.100 300.000 138.300 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 141.180 300.000 142.380 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 145.260 300.000 146.460 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 148.660 300.000 149.860 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 152.740 300.000 153.940 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 156.140 300.000 157.340 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.030 296.000 229.590 300.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.610 0.000 56.170 4.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 270.380 300.000 271.580 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.330 0.000 93.890 4.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.590 0.000 131.150 4.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.310 0.000 168.870 4.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 280.580 4.000 281.780 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 273.780 300.000 274.980 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.570 0.000 206.130 4.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.090 296.000 257.650 300.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 277.860 300.000 279.060 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.550 296.000 235.110 300.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.290 0.000 243.850 4.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.610 296.000 263.170 300.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.590 296.000 269.150 300.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.110 296.000 274.670 300.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.660 4.000 285.860 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 281.940 300.000 283.140 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.630 296.000 280.190 300.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 285.340 300.000 286.540 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 288.740 4.000 289.940 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 289.420 300.000 290.620 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.070 296.000 240.630 300.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.550 0.000 281.110 4.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.610 296.000 286.170 300.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.130 296.000 291.690 300.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.820 4.000 294.020 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 292.820 300.000 294.020 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 296.900 4.000 298.100 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 296.900 300.000 298.100 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.650 296.000 297.210 300.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.350 0.000 18.910 4.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 268.340 4.000 269.540 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 266.300 300.000 267.500 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.420 4.000 273.620 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.590 296.000 246.150 300.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.570 296.000 252.130 300.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 276.500 4.000 277.700 ;
    END
  END io_out[9]
  PIN la1_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1.780 4.000 2.980 ;
    END
  END la1_data_in[0]
  PIN la1_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.260 4.000 44.460 ;
    END
  END la1_data_in[10]
  PIN la1_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.340 4.000 48.540 ;
    END
  END la1_data_in[11]
  PIN la1_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.420 4.000 52.620 ;
    END
  END la1_data_in[12]
  PIN la1_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.500 4.000 56.700 ;
    END
  END la1_data_in[13]
  PIN la1_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.580 4.000 60.780 ;
    END
  END la1_data_in[14]
  PIN la1_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.660 4.000 64.860 ;
    END
  END la1_data_in[15]
  PIN la1_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.420 4.000 69.620 ;
    END
  END la1_data_in[16]
  PIN la1_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.500 4.000 73.700 ;
    END
  END la1_data_in[17]
  PIN la1_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.580 4.000 77.780 ;
    END
  END la1_data_in[18]
  PIN la1_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.660 4.000 81.860 ;
    END
  END la1_data_in[19]
  PIN la1_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 5.860 4.000 7.060 ;
    END
  END la1_data_in[1]
  PIN la1_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.740 4.000 85.940 ;
    END
  END la1_data_in[20]
  PIN la1_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.820 4.000 90.020 ;
    END
  END la1_data_in[21]
  PIN la1_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.900 4.000 94.100 ;
    END
  END la1_data_in[22]
  PIN la1_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.980 4.000 98.180 ;
    END
  END la1_data_in[23]
  PIN la1_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 101.740 4.000 102.940 ;
    END
  END la1_data_in[24]
  PIN la1_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.820 4.000 107.020 ;
    END
  END la1_data_in[25]
  PIN la1_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 109.900 4.000 111.100 ;
    END
  END la1_data_in[26]
  PIN la1_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 113.980 4.000 115.180 ;
    END
  END la1_data_in[27]
  PIN la1_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.060 4.000 119.260 ;
    END
  END la1_data_in[28]
  PIN la1_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.140 4.000 123.340 ;
    END
  END la1_data_in[29]
  PIN la1_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 9.940 4.000 11.140 ;
    END
  END la1_data_in[2]
  PIN la1_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.220 4.000 127.420 ;
    END
  END la1_data_in[30]
  PIN la1_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.300 4.000 131.500 ;
    END
  END la1_data_in[31]
  PIN la1_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 14.020 4.000 15.220 ;
    END
  END la1_data_in[3]
  PIN la1_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 18.100 4.000 19.300 ;
    END
  END la1_data_in[4]
  PIN la1_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 22.180 4.000 23.380 ;
    END
  END la1_data_in[5]
  PIN la1_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 26.260 4.000 27.460 ;
    END
  END la1_data_in[6]
  PIN la1_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.340 4.000 31.540 ;
    END
  END la1_data_in[7]
  PIN la1_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.100 4.000 36.300 ;
    END
  END la1_data_in[8]
  PIN la1_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.180 4.000 40.380 ;
    END
  END la1_data_in[9]
  PIN la1_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 135.060 4.000 136.260 ;
    END
  END la1_data_out[0]
  PIN la1_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.540 4.000 177.740 ;
    END
  END la1_data_out[10]
  PIN la1_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.620 4.000 181.820 ;
    END
  END la1_data_out[11]
  PIN la1_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 184.700 4.000 185.900 ;
    END
  END la1_data_out[12]
  PIN la1_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 188.780 4.000 189.980 ;
    END
  END la1_data_out[13]
  PIN la1_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 192.860 4.000 194.060 ;
    END
  END la1_data_out[14]
  PIN la1_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 196.940 4.000 198.140 ;
    END
  END la1_data_out[15]
  PIN la1_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 201.700 4.000 202.900 ;
    END
  END la1_data_out[16]
  PIN la1_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 205.780 4.000 206.980 ;
    END
  END la1_data_out[17]
  PIN la1_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.860 4.000 211.060 ;
    END
  END la1_data_out[18]
  PIN la1_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 213.940 4.000 215.140 ;
    END
  END la1_data_out[19]
  PIN la1_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.140 4.000 140.340 ;
    END
  END la1_data_out[1]
  PIN la1_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 218.020 4.000 219.220 ;
    END
  END la1_data_out[20]
  PIN la1_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 222.100 4.000 223.300 ;
    END
  END la1_data_out[21]
  PIN la1_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 226.180 4.000 227.380 ;
    END
  END la1_data_out[22]
  PIN la1_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 230.260 4.000 231.460 ;
    END
  END la1_data_out[23]
  PIN la1_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 235.020 4.000 236.220 ;
    END
  END la1_data_out[24]
  PIN la1_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 239.100 4.000 240.300 ;
    END
  END la1_data_out[25]
  PIN la1_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 243.180 4.000 244.380 ;
    END
  END la1_data_out[26]
  PIN la1_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 247.260 4.000 248.460 ;
    END
  END la1_data_out[27]
  PIN la1_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.340 4.000 252.540 ;
    END
  END la1_data_out[28]
  PIN la1_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.420 4.000 256.620 ;
    END
  END la1_data_out[29]
  PIN la1_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 143.220 4.000 144.420 ;
    END
  END la1_data_out[2]
  PIN la1_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.500 4.000 260.700 ;
    END
  END la1_data_out[30]
  PIN la1_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 263.580 4.000 264.780 ;
    END
  END la1_data_out[31]
  PIN la1_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 147.300 4.000 148.500 ;
    END
  END la1_data_out[3]
  PIN la1_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.380 4.000 152.580 ;
    END
  END la1_data_out[4]
  PIN la1_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.460 4.000 156.660 ;
    END
  END la1_data_out[5]
  PIN la1_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.540 4.000 160.740 ;
    END
  END la1_data_out[6]
  PIN la1_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.620 4.000 164.820 ;
    END
  END la1_data_out[7]
  PIN la1_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.380 4.000 169.580 ;
    END
  END la1_data_out[8]
  PIN la1_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.460 4.000 173.660 ;
    END
  END la1_data_out[9]
  PIN la1_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 1.100 300.000 2.300 ;
    END
  END la1_oenb[0]
  PIN la1_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 38.500 300.000 39.700 ;
    END
  END la1_oenb[10]
  PIN la1_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 42.580 300.000 43.780 ;
    END
  END la1_oenb[11]
  PIN la1_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 45.980 300.000 47.180 ;
    END
  END la1_oenb[12]
  PIN la1_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 50.060 300.000 51.260 ;
    END
  END la1_oenb[13]
  PIN la1_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 54.140 300.000 55.340 ;
    END
  END la1_oenb[14]
  PIN la1_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 57.540 300.000 58.740 ;
    END
  END la1_oenb[15]
  PIN la1_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 61.620 300.000 62.820 ;
    END
  END la1_oenb[16]
  PIN la1_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 65.020 300.000 66.220 ;
    END
  END la1_oenb[17]
  PIN la1_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 69.100 300.000 70.300 ;
    END
  END la1_oenb[18]
  PIN la1_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 73.180 300.000 74.380 ;
    END
  END la1_oenb[19]
  PIN la1_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 4.500 300.000 5.700 ;
    END
  END la1_oenb[1]
  PIN la1_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 76.580 300.000 77.780 ;
    END
  END la1_oenb[20]
  PIN la1_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 80.660 300.000 81.860 ;
    END
  END la1_oenb[21]
  PIN la1_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 84.060 300.000 85.260 ;
    END
  END la1_oenb[22]
  PIN la1_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 88.140 300.000 89.340 ;
    END
  END la1_oenb[23]
  PIN la1_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 91.540 300.000 92.740 ;
    END
  END la1_oenb[24]
  PIN la1_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 95.620 300.000 96.820 ;
    END
  END la1_oenb[25]
  PIN la1_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 99.700 300.000 100.900 ;
    END
  END la1_oenb[26]
  PIN la1_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 103.100 300.000 104.300 ;
    END
  END la1_oenb[27]
  PIN la1_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 107.180 300.000 108.380 ;
    END
  END la1_oenb[28]
  PIN la1_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 110.580 300.000 111.780 ;
    END
  END la1_oenb[29]
  PIN la1_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 8.580 300.000 9.780 ;
    END
  END la1_oenb[2]
  PIN la1_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 114.660 300.000 115.860 ;
    END
  END la1_oenb[30]
  PIN la1_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 118.740 300.000 119.940 ;
    END
  END la1_oenb[31]
  PIN la1_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 11.980 300.000 13.180 ;
    END
  END la1_oenb[3]
  PIN la1_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 16.060 300.000 17.260 ;
    END
  END la1_oenb[4]
  PIN la1_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 19.460 300.000 20.660 ;
    END
  END la1_oenb[5]
  PIN la1_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 23.540 300.000 24.740 ;
    END
  END la1_oenb[6]
  PIN la1_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 27.620 300.000 28.820 ;
    END
  END la1_oenb[7]
  PIN la1_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 31.020 300.000 32.220 ;
    END
  END la1_oenb[8]
  PIN la1_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 35.100 300.000 36.300 ;
    END
  END la1_oenb[9]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 2.480 22.640 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 2.480 176.240 288.560 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 2.480 99.440 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 2.480 253.040 288.560 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.230 296.000 8.790 300.000 ;
    END
  END wb_clk_i
  OBS
      LAYER li1 ;
        RECT 5.520 2.635 294.400 288.405 ;
      LAYER met1 ;
        RECT 2.830 1.400 297.090 288.960 ;
      LAYER met2 ;
        RECT 3.550 295.720 7.950 297.685 ;
        RECT 9.070 295.720 13.470 297.685 ;
        RECT 14.590 295.720 18.990 297.685 ;
        RECT 20.110 295.720 24.970 297.685 ;
        RECT 26.090 295.720 30.490 297.685 ;
        RECT 31.610 295.720 36.010 297.685 ;
        RECT 37.130 295.720 41.990 297.685 ;
        RECT 43.110 295.720 47.510 297.685 ;
        RECT 48.630 295.720 53.030 297.685 ;
        RECT 54.150 295.720 59.010 297.685 ;
        RECT 60.130 295.720 64.530 297.685 ;
        RECT 65.650 295.720 70.050 297.685 ;
        RECT 71.170 295.720 75.570 297.685 ;
        RECT 76.690 295.720 81.550 297.685 ;
        RECT 82.670 295.720 87.070 297.685 ;
        RECT 88.190 295.720 92.590 297.685 ;
        RECT 93.710 295.720 98.570 297.685 ;
        RECT 99.690 295.720 104.090 297.685 ;
        RECT 105.210 295.720 109.610 297.685 ;
        RECT 110.730 295.720 115.590 297.685 ;
        RECT 116.710 295.720 121.110 297.685 ;
        RECT 122.230 295.720 126.630 297.685 ;
        RECT 127.750 295.720 132.150 297.685 ;
        RECT 133.270 295.720 138.130 297.685 ;
        RECT 139.250 295.720 143.650 297.685 ;
        RECT 144.770 295.720 149.170 297.685 ;
        RECT 150.290 295.720 155.150 297.685 ;
        RECT 156.270 295.720 160.670 297.685 ;
        RECT 161.790 295.720 166.190 297.685 ;
        RECT 167.310 295.720 172.170 297.685 ;
        RECT 173.290 295.720 177.690 297.685 ;
        RECT 178.810 295.720 183.210 297.685 ;
        RECT 184.330 295.720 188.730 297.685 ;
        RECT 189.850 295.720 194.710 297.685 ;
        RECT 195.830 295.720 200.230 297.685 ;
        RECT 201.350 295.720 205.750 297.685 ;
        RECT 206.870 295.720 211.730 297.685 ;
        RECT 212.850 295.720 217.250 297.685 ;
        RECT 218.370 295.720 222.770 297.685 ;
        RECT 223.890 295.720 228.750 297.685 ;
        RECT 229.870 295.720 234.270 297.685 ;
        RECT 235.390 295.720 239.790 297.685 ;
        RECT 240.910 295.720 245.310 297.685 ;
        RECT 246.430 295.720 251.290 297.685 ;
        RECT 252.410 295.720 256.810 297.685 ;
        RECT 257.930 295.720 262.330 297.685 ;
        RECT 263.450 295.720 268.310 297.685 ;
        RECT 269.430 295.720 273.830 297.685 ;
        RECT 274.950 295.720 279.350 297.685 ;
        RECT 280.470 295.720 285.330 297.685 ;
        RECT 286.450 295.720 290.850 297.685 ;
        RECT 291.970 295.720 296.370 297.685 ;
        RECT 2.860 4.280 297.060 295.720 ;
        RECT 2.860 1.370 18.070 4.280 ;
        RECT 19.190 1.370 55.330 4.280 ;
        RECT 56.450 1.370 93.050 4.280 ;
        RECT 94.170 1.370 130.310 4.280 ;
        RECT 131.430 1.370 168.030 4.280 ;
        RECT 169.150 1.370 205.290 4.280 ;
        RECT 206.410 1.370 243.010 4.280 ;
        RECT 244.130 1.370 280.270 4.280 ;
        RECT 281.390 1.370 297.060 4.280 ;
      LAYER met3 ;
        RECT 4.400 296.500 295.600 297.665 ;
        RECT 4.000 294.420 296.000 296.500 ;
        RECT 4.400 292.420 295.600 294.420 ;
        RECT 4.000 291.020 296.000 292.420 ;
        RECT 4.000 290.340 295.600 291.020 ;
        RECT 4.400 289.020 295.600 290.340 ;
        RECT 4.400 288.340 296.000 289.020 ;
        RECT 4.000 286.940 296.000 288.340 ;
        RECT 4.000 286.260 295.600 286.940 ;
        RECT 4.400 284.940 295.600 286.260 ;
        RECT 4.400 284.260 296.000 284.940 ;
        RECT 4.000 283.540 296.000 284.260 ;
        RECT 4.000 282.180 295.600 283.540 ;
        RECT 4.400 281.540 295.600 282.180 ;
        RECT 4.400 280.180 296.000 281.540 ;
        RECT 4.000 279.460 296.000 280.180 ;
        RECT 4.000 278.100 295.600 279.460 ;
        RECT 4.400 277.460 295.600 278.100 ;
        RECT 4.400 276.100 296.000 277.460 ;
        RECT 4.000 275.380 296.000 276.100 ;
        RECT 4.000 274.020 295.600 275.380 ;
        RECT 4.400 273.380 295.600 274.020 ;
        RECT 4.400 272.020 296.000 273.380 ;
        RECT 4.000 271.980 296.000 272.020 ;
        RECT 4.000 269.980 295.600 271.980 ;
        RECT 4.000 269.940 296.000 269.980 ;
        RECT 4.400 267.940 296.000 269.940 ;
        RECT 4.000 267.900 296.000 267.940 ;
        RECT 4.000 265.900 295.600 267.900 ;
        RECT 4.000 265.180 296.000 265.900 ;
        RECT 4.400 264.500 296.000 265.180 ;
        RECT 4.400 263.180 295.600 264.500 ;
        RECT 4.000 262.500 295.600 263.180 ;
        RECT 4.000 261.100 296.000 262.500 ;
        RECT 4.400 260.420 296.000 261.100 ;
        RECT 4.400 259.100 295.600 260.420 ;
        RECT 4.000 258.420 295.600 259.100 ;
        RECT 4.000 257.020 296.000 258.420 ;
        RECT 4.400 255.020 295.600 257.020 ;
        RECT 4.000 252.940 296.000 255.020 ;
        RECT 4.400 250.940 295.600 252.940 ;
        RECT 4.000 248.860 296.000 250.940 ;
        RECT 4.400 246.860 295.600 248.860 ;
        RECT 4.000 245.460 296.000 246.860 ;
        RECT 4.000 244.780 295.600 245.460 ;
        RECT 4.400 243.460 295.600 244.780 ;
        RECT 4.400 242.780 296.000 243.460 ;
        RECT 4.000 241.380 296.000 242.780 ;
        RECT 4.000 240.700 295.600 241.380 ;
        RECT 4.400 239.380 295.600 240.700 ;
        RECT 4.400 238.700 296.000 239.380 ;
        RECT 4.000 237.980 296.000 238.700 ;
        RECT 4.000 236.620 295.600 237.980 ;
        RECT 4.400 235.980 295.600 236.620 ;
        RECT 4.400 234.620 296.000 235.980 ;
        RECT 4.000 233.900 296.000 234.620 ;
        RECT 4.000 231.900 295.600 233.900 ;
        RECT 4.000 231.860 296.000 231.900 ;
        RECT 4.400 229.860 296.000 231.860 ;
        RECT 4.000 229.820 296.000 229.860 ;
        RECT 4.000 227.820 295.600 229.820 ;
        RECT 4.000 227.780 296.000 227.820 ;
        RECT 4.400 226.420 296.000 227.780 ;
        RECT 4.400 225.780 295.600 226.420 ;
        RECT 4.000 224.420 295.600 225.780 ;
        RECT 4.000 223.700 296.000 224.420 ;
        RECT 4.400 222.340 296.000 223.700 ;
        RECT 4.400 221.700 295.600 222.340 ;
        RECT 4.000 220.340 295.600 221.700 ;
        RECT 4.000 219.620 296.000 220.340 ;
        RECT 4.400 218.940 296.000 219.620 ;
        RECT 4.400 217.620 295.600 218.940 ;
        RECT 4.000 216.940 295.600 217.620 ;
        RECT 4.000 215.540 296.000 216.940 ;
        RECT 4.400 214.860 296.000 215.540 ;
        RECT 4.400 213.540 295.600 214.860 ;
        RECT 4.000 212.860 295.600 213.540 ;
        RECT 4.000 211.460 296.000 212.860 ;
        RECT 4.400 209.460 295.600 211.460 ;
        RECT 4.000 207.380 296.000 209.460 ;
        RECT 4.400 205.380 295.600 207.380 ;
        RECT 4.000 203.300 296.000 205.380 ;
        RECT 4.400 201.300 295.600 203.300 ;
        RECT 4.000 199.900 296.000 201.300 ;
        RECT 4.000 198.540 295.600 199.900 ;
        RECT 4.400 197.900 295.600 198.540 ;
        RECT 4.400 196.540 296.000 197.900 ;
        RECT 4.000 195.820 296.000 196.540 ;
        RECT 4.000 194.460 295.600 195.820 ;
        RECT 4.400 193.820 295.600 194.460 ;
        RECT 4.400 192.460 296.000 193.820 ;
        RECT 4.000 192.420 296.000 192.460 ;
        RECT 4.000 190.420 295.600 192.420 ;
        RECT 4.000 190.380 296.000 190.420 ;
        RECT 4.400 188.380 296.000 190.380 ;
        RECT 4.000 188.340 296.000 188.380 ;
        RECT 4.000 186.340 295.600 188.340 ;
        RECT 4.000 186.300 296.000 186.340 ;
        RECT 4.400 184.300 296.000 186.300 ;
        RECT 4.000 184.260 296.000 184.300 ;
        RECT 4.000 182.260 295.600 184.260 ;
        RECT 4.000 182.220 296.000 182.260 ;
        RECT 4.400 180.860 296.000 182.220 ;
        RECT 4.400 180.220 295.600 180.860 ;
        RECT 4.000 178.860 295.600 180.220 ;
        RECT 4.000 178.140 296.000 178.860 ;
        RECT 4.400 176.780 296.000 178.140 ;
        RECT 4.400 176.140 295.600 176.780 ;
        RECT 4.000 174.780 295.600 176.140 ;
        RECT 4.000 174.060 296.000 174.780 ;
        RECT 4.400 173.380 296.000 174.060 ;
        RECT 4.400 172.060 295.600 173.380 ;
        RECT 4.000 171.380 295.600 172.060 ;
        RECT 4.000 169.980 296.000 171.380 ;
        RECT 4.400 169.300 296.000 169.980 ;
        RECT 4.400 167.980 295.600 169.300 ;
        RECT 4.000 167.300 295.600 167.980 ;
        RECT 4.000 165.900 296.000 167.300 ;
        RECT 4.000 165.220 295.600 165.900 ;
        RECT 4.400 163.900 295.600 165.220 ;
        RECT 4.400 163.220 296.000 163.900 ;
        RECT 4.000 161.820 296.000 163.220 ;
        RECT 4.000 161.140 295.600 161.820 ;
        RECT 4.400 159.820 295.600 161.140 ;
        RECT 4.400 159.140 296.000 159.820 ;
        RECT 4.000 157.740 296.000 159.140 ;
        RECT 4.000 157.060 295.600 157.740 ;
        RECT 4.400 155.740 295.600 157.060 ;
        RECT 4.400 155.060 296.000 155.740 ;
        RECT 4.000 154.340 296.000 155.060 ;
        RECT 4.000 152.980 295.600 154.340 ;
        RECT 4.400 152.340 295.600 152.980 ;
        RECT 4.400 150.980 296.000 152.340 ;
        RECT 4.000 150.260 296.000 150.980 ;
        RECT 4.000 148.900 295.600 150.260 ;
        RECT 4.400 148.260 295.600 148.900 ;
        RECT 4.400 146.900 296.000 148.260 ;
        RECT 4.000 146.860 296.000 146.900 ;
        RECT 4.000 144.860 295.600 146.860 ;
        RECT 4.000 144.820 296.000 144.860 ;
        RECT 4.400 142.820 296.000 144.820 ;
        RECT 4.000 142.780 296.000 142.820 ;
        RECT 4.000 140.780 295.600 142.780 ;
        RECT 4.000 140.740 296.000 140.780 ;
        RECT 4.400 138.740 296.000 140.740 ;
        RECT 4.000 138.700 296.000 138.740 ;
        RECT 4.000 136.700 295.600 138.700 ;
        RECT 4.000 136.660 296.000 136.700 ;
        RECT 4.400 135.300 296.000 136.660 ;
        RECT 4.400 134.660 295.600 135.300 ;
        RECT 4.000 133.300 295.600 134.660 ;
        RECT 4.000 131.900 296.000 133.300 ;
        RECT 4.400 131.220 296.000 131.900 ;
        RECT 4.400 129.900 295.600 131.220 ;
        RECT 4.000 129.220 295.600 129.900 ;
        RECT 4.000 127.820 296.000 129.220 ;
        RECT 4.400 125.820 295.600 127.820 ;
        RECT 4.000 123.740 296.000 125.820 ;
        RECT 4.400 121.740 295.600 123.740 ;
        RECT 4.000 120.340 296.000 121.740 ;
        RECT 4.000 119.660 295.600 120.340 ;
        RECT 4.400 118.340 295.600 119.660 ;
        RECT 4.400 117.660 296.000 118.340 ;
        RECT 4.000 116.260 296.000 117.660 ;
        RECT 4.000 115.580 295.600 116.260 ;
        RECT 4.400 114.260 295.600 115.580 ;
        RECT 4.400 113.580 296.000 114.260 ;
        RECT 4.000 112.180 296.000 113.580 ;
        RECT 4.000 111.500 295.600 112.180 ;
        RECT 4.400 110.180 295.600 111.500 ;
        RECT 4.400 109.500 296.000 110.180 ;
        RECT 4.000 108.780 296.000 109.500 ;
        RECT 4.000 107.420 295.600 108.780 ;
        RECT 4.400 106.780 295.600 107.420 ;
        RECT 4.400 105.420 296.000 106.780 ;
        RECT 4.000 104.700 296.000 105.420 ;
        RECT 4.000 103.340 295.600 104.700 ;
        RECT 4.400 102.700 295.600 103.340 ;
        RECT 4.400 101.340 296.000 102.700 ;
        RECT 4.000 101.300 296.000 101.340 ;
        RECT 4.000 99.300 295.600 101.300 ;
        RECT 4.000 98.580 296.000 99.300 ;
        RECT 4.400 97.220 296.000 98.580 ;
        RECT 4.400 96.580 295.600 97.220 ;
        RECT 4.000 95.220 295.600 96.580 ;
        RECT 4.000 94.500 296.000 95.220 ;
        RECT 4.400 93.140 296.000 94.500 ;
        RECT 4.400 92.500 295.600 93.140 ;
        RECT 4.000 91.140 295.600 92.500 ;
        RECT 4.000 90.420 296.000 91.140 ;
        RECT 4.400 89.740 296.000 90.420 ;
        RECT 4.400 88.420 295.600 89.740 ;
        RECT 4.000 87.740 295.600 88.420 ;
        RECT 4.000 86.340 296.000 87.740 ;
        RECT 4.400 85.660 296.000 86.340 ;
        RECT 4.400 84.340 295.600 85.660 ;
        RECT 4.000 83.660 295.600 84.340 ;
        RECT 4.000 82.260 296.000 83.660 ;
        RECT 4.400 80.260 295.600 82.260 ;
        RECT 4.000 78.180 296.000 80.260 ;
        RECT 4.400 76.180 295.600 78.180 ;
        RECT 4.000 74.780 296.000 76.180 ;
        RECT 4.000 74.100 295.600 74.780 ;
        RECT 4.400 72.780 295.600 74.100 ;
        RECT 4.400 72.100 296.000 72.780 ;
        RECT 4.000 70.700 296.000 72.100 ;
        RECT 4.000 70.020 295.600 70.700 ;
        RECT 4.400 68.700 295.600 70.020 ;
        RECT 4.400 68.020 296.000 68.700 ;
        RECT 4.000 66.620 296.000 68.020 ;
        RECT 4.000 65.260 295.600 66.620 ;
        RECT 4.400 64.620 295.600 65.260 ;
        RECT 4.400 63.260 296.000 64.620 ;
        RECT 4.000 63.220 296.000 63.260 ;
        RECT 4.000 61.220 295.600 63.220 ;
        RECT 4.000 61.180 296.000 61.220 ;
        RECT 4.400 59.180 296.000 61.180 ;
        RECT 4.000 59.140 296.000 59.180 ;
        RECT 4.000 57.140 295.600 59.140 ;
        RECT 4.000 57.100 296.000 57.140 ;
        RECT 4.400 55.740 296.000 57.100 ;
        RECT 4.400 55.100 295.600 55.740 ;
        RECT 4.000 53.740 295.600 55.100 ;
        RECT 4.000 53.020 296.000 53.740 ;
        RECT 4.400 51.660 296.000 53.020 ;
        RECT 4.400 51.020 295.600 51.660 ;
        RECT 4.000 49.660 295.600 51.020 ;
        RECT 4.000 48.940 296.000 49.660 ;
        RECT 4.400 47.580 296.000 48.940 ;
        RECT 4.400 46.940 295.600 47.580 ;
        RECT 4.000 45.580 295.600 46.940 ;
        RECT 4.000 44.860 296.000 45.580 ;
        RECT 4.400 44.180 296.000 44.860 ;
        RECT 4.400 42.860 295.600 44.180 ;
        RECT 4.000 42.180 295.600 42.860 ;
        RECT 4.000 40.780 296.000 42.180 ;
        RECT 4.400 40.100 296.000 40.780 ;
        RECT 4.400 38.780 295.600 40.100 ;
        RECT 4.000 38.100 295.600 38.780 ;
        RECT 4.000 36.700 296.000 38.100 ;
        RECT 4.400 34.700 295.600 36.700 ;
        RECT 4.000 32.620 296.000 34.700 ;
        RECT 4.000 31.940 295.600 32.620 ;
        RECT 4.400 30.620 295.600 31.940 ;
        RECT 4.400 29.940 296.000 30.620 ;
        RECT 4.000 29.220 296.000 29.940 ;
        RECT 4.000 27.860 295.600 29.220 ;
        RECT 4.400 27.220 295.600 27.860 ;
        RECT 4.400 25.860 296.000 27.220 ;
        RECT 4.000 25.140 296.000 25.860 ;
        RECT 4.000 23.780 295.600 25.140 ;
        RECT 4.400 23.140 295.600 23.780 ;
        RECT 4.400 21.780 296.000 23.140 ;
        RECT 4.000 21.060 296.000 21.780 ;
        RECT 4.000 19.700 295.600 21.060 ;
        RECT 4.400 19.060 295.600 19.700 ;
        RECT 4.400 17.700 296.000 19.060 ;
        RECT 4.000 17.660 296.000 17.700 ;
        RECT 4.000 15.660 295.600 17.660 ;
        RECT 4.000 15.620 296.000 15.660 ;
        RECT 4.400 13.620 296.000 15.620 ;
        RECT 4.000 13.580 296.000 13.620 ;
        RECT 4.000 11.580 295.600 13.580 ;
        RECT 4.000 11.540 296.000 11.580 ;
        RECT 4.400 10.180 296.000 11.540 ;
        RECT 4.400 9.540 295.600 10.180 ;
        RECT 4.000 8.180 295.600 9.540 ;
        RECT 4.000 7.460 296.000 8.180 ;
        RECT 4.400 6.100 296.000 7.460 ;
        RECT 4.400 5.460 295.600 6.100 ;
        RECT 4.000 4.100 295.600 5.460 ;
        RECT 4.000 3.380 296.000 4.100 ;
        RECT 4.400 2.700 296.000 3.380 ;
        RECT 4.400 2.555 295.600 2.700 ;
      LAYER met4 ;
        RECT 62.855 6.295 97.440 283.385 ;
        RECT 99.840 6.295 174.240 283.385 ;
        RECT 176.640 6.295 228.785 283.385 ;
  END
END wrapped_vgademo_on_fpga
END LIBRARY

