VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_vgademo_on_fpga
  CLASS BLOCK ;
  FOREIGN wrapped_vgademo_on_fpga ;
  ORIGIN 0.000 0.000 ;
  SIZE 300.000 BY 300.000 ;
  PIN active
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.170 296.000 3.730 300.000 ;
    END
  END active
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.050 296.000 16.610 300.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.370 296.000 81.930 300.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.810 296.000 88.370 300.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.250 296.000 94.810 300.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.690 296.000 101.250 300.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.130 296.000 107.690 300.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.570 296.000 114.130 300.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.470 296.000 121.030 300.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.910 296.000 127.470 300.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.350 296.000 133.910 300.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.790 296.000 140.350 300.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.490 296.000 23.050 300.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.230 296.000 146.790 300.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.130 296.000 153.690 300.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.570 296.000 160.130 300.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.010 296.000 166.570 300.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.450 296.000 173.010 300.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.890 296.000 179.450 300.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.330 296.000 185.890 300.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.230 296.000 192.790 300.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.670 296.000 199.230 300.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.110 296.000 205.670 300.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.930 296.000 29.490 300.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.550 296.000 212.110 300.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.990 296.000 218.550 300.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.430 296.000 224.990 300.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.330 296.000 231.890 300.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.770 296.000 238.330 300.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.210 296.000 244.770 300.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.650 296.000 251.210 300.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.090 296.000 257.650 300.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.370 296.000 35.930 300.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.270 296.000 42.830 300.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.710 296.000 49.270 300.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.150 296.000 55.710 300.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.590 296.000 62.150 300.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.030 296.000 68.590 300.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.470 296.000 75.030 300.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 120.780 300.000 121.980 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 158.180 300.000 159.380 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 162.260 300.000 163.460 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 165.660 300.000 166.860 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 169.740 300.000 170.940 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 173.140 300.000 174.340 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 177.220 300.000 178.420 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 180.620 300.000 181.820 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 184.700 300.000 185.900 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 188.100 300.000 189.300 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 192.180 300.000 193.380 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 124.180 300.000 125.380 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 195.580 300.000 196.780 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 199.660 300.000 200.860 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 203.060 300.000 204.260 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 207.140 300.000 208.340 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 210.540 300.000 211.740 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 214.620 300.000 215.820 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 218.020 300.000 219.220 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 222.100 300.000 223.300 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 225.500 300.000 226.700 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 229.580 300.000 230.780 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 128.260 300.000 129.460 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 232.980 300.000 234.180 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 237.060 300.000 238.260 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 240.460 300.000 241.660 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 244.540 300.000 245.740 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 247.940 300.000 249.140 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 252.020 300.000 253.220 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 255.420 300.000 256.620 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 259.500 300.000 260.700 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 131.660 300.000 132.860 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 135.740 300.000 136.940 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 139.140 300.000 140.340 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 143.220 300.000 144.420 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 146.620 300.000 147.820 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 150.700 300.000 151.900 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 154.780 300.000 155.980 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 256.780 4.000 257.980 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 270.380 300.000 271.580 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.710 0.000 95.270 4.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.870 296.000 277.430 300.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 268.340 4.000 269.540 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.310 0.000 122.870 4.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 274.460 300.000 275.660 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.450 0.000 150.010 4.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.590 0.000 177.150 4.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.730 0.000 204.290 4.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.330 0.000 231.890 4.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.290 0.000 13.850 4.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.420 4.000 273.620 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.470 0.000 259.030 4.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 276.500 4.000 277.700 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 277.860 300.000 279.060 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.610 0.000 286.170 4.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 280.580 4.000 281.780 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.660 4.000 285.860 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 281.940 300.000 283.140 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 288.740 4.000 289.940 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 285.340 300.000 286.540 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 262.900 300.000 264.100 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.310 296.000 283.870 300.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 289.420 300.000 290.620 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.820 4.000 294.020 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 296.900 4.000 298.100 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.750 296.000 290.310 300.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 292.820 300.000 294.020 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 296.900 300.000 298.100 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.190 296.000 296.750 300.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.530 296.000 264.090 300.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 260.860 4.000 262.060 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 264.940 4.000 266.140 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.430 296.000 270.990 300.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 266.980 300.000 268.180 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.430 0.000 40.990 4.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.570 0.000 68.130 4.000 ;
    END
  END io_out[9]
  PIN la1_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1.100 4.000 2.300 ;
    END
  END la1_data_in[0]
  PIN la1_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.540 4.000 41.740 ;
    END
  END la1_data_in[10]
  PIN la1_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.620 4.000 45.820 ;
    END
  END la1_data_in[11]
  PIN la1_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.700 4.000 49.900 ;
    END
  END la1_data_in[12]
  PIN la1_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 52.780 4.000 53.980 ;
    END
  END la1_data_in[13]
  PIN la1_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 56.860 4.000 58.060 ;
    END
  END la1_data_in[14]
  PIN la1_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 60.940 4.000 62.140 ;
    END
  END la1_data_in[15]
  PIN la1_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.020 4.000 66.220 ;
    END
  END la1_data_in[16]
  PIN la1_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.420 4.000 69.620 ;
    END
  END la1_data_in[17]
  PIN la1_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.500 4.000 73.700 ;
    END
  END la1_data_in[18]
  PIN la1_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.580 4.000 77.780 ;
    END
  END la1_data_in[19]
  PIN la1_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.500 4.000 5.700 ;
    END
  END la1_data_in[1]
  PIN la1_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.660 4.000 81.860 ;
    END
  END la1_data_in[20]
  PIN la1_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.740 4.000 85.940 ;
    END
  END la1_data_in[21]
  PIN la1_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.820 4.000 90.020 ;
    END
  END la1_data_in[22]
  PIN la1_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.900 4.000 94.100 ;
    END
  END la1_data_in[23]
  PIN la1_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.980 4.000 98.180 ;
    END
  END la1_data_in[24]
  PIN la1_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 101.060 4.000 102.260 ;
    END
  END la1_data_in[25]
  PIN la1_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.460 4.000 105.660 ;
    END
  END la1_data_in[26]
  PIN la1_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.540 4.000 109.740 ;
    END
  END la1_data_in[27]
  PIN la1_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.620 4.000 113.820 ;
    END
  END la1_data_in[28]
  PIN la1_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 116.700 4.000 117.900 ;
    END
  END la1_data_in[29]
  PIN la1_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.580 4.000 9.780 ;
    END
  END la1_data_in[2]
  PIN la1_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 120.780 4.000 121.980 ;
    END
  END la1_data_in[30]
  PIN la1_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 124.860 4.000 126.060 ;
    END
  END la1_data_in[31]
  PIN la1_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.660 4.000 13.860 ;
    END
  END la1_data_in[3]
  PIN la1_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.740 4.000 17.940 ;
    END
  END la1_data_in[4]
  PIN la1_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.820 4.000 22.020 ;
    END
  END la1_data_in[5]
  PIN la1_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.900 4.000 26.100 ;
    END
  END la1_data_in[6]
  PIN la1_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.980 4.000 30.180 ;
    END
  END la1_data_in[7]
  PIN la1_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.060 4.000 34.260 ;
    END
  END la1_data_in[8]
  PIN la1_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.460 4.000 37.660 ;
    END
  END la1_data_in[9]
  PIN la1_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 128.940 4.000 130.140 ;
    END
  END la1_data_out[0]
  PIN la1_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.380 4.000 169.580 ;
    END
  END la1_data_out[10]
  PIN la1_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.460 4.000 173.660 ;
    END
  END la1_data_out[11]
  PIN la1_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.540 4.000 177.740 ;
    END
  END la1_data_out[12]
  PIN la1_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.620 4.000 181.820 ;
    END
  END la1_data_out[13]
  PIN la1_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 184.700 4.000 185.900 ;
    END
  END la1_data_out[14]
  PIN la1_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 188.780 4.000 189.980 ;
    END
  END la1_data_out[15]
  PIN la1_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 192.860 4.000 194.060 ;
    END
  END la1_data_out[16]
  PIN la1_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 196.940 4.000 198.140 ;
    END
  END la1_data_out[17]
  PIN la1_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 201.020 4.000 202.220 ;
    END
  END la1_data_out[18]
  PIN la1_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.420 4.000 205.620 ;
    END
  END la1_data_out[19]
  PIN la1_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 133.020 4.000 134.220 ;
    END
  END la1_data_out[1]
  PIN la1_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.500 4.000 209.700 ;
    END
  END la1_data_out[20]
  PIN la1_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.580 4.000 213.780 ;
    END
  END la1_data_out[21]
  PIN la1_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.660 4.000 217.860 ;
    END
  END la1_data_out[22]
  PIN la1_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 220.740 4.000 221.940 ;
    END
  END la1_data_out[23]
  PIN la1_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.820 4.000 226.020 ;
    END
  END la1_data_out[24]
  PIN la1_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 228.900 4.000 230.100 ;
    END
  END la1_data_out[25]
  PIN la1_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 232.980 4.000 234.180 ;
    END
  END la1_data_out[26]
  PIN la1_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.380 4.000 237.580 ;
    END
  END la1_data_out[27]
  PIN la1_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.460 4.000 241.660 ;
    END
  END la1_data_out[28]
  PIN la1_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.540 4.000 245.740 ;
    END
  END la1_data_out[29]
  PIN la1_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.420 4.000 137.620 ;
    END
  END la1_data_out[2]
  PIN la1_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.620 4.000 249.820 ;
    END
  END la1_data_out[30]
  PIN la1_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 252.700 4.000 253.900 ;
    END
  END la1_data_out[31]
  PIN la1_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.500 4.000 141.700 ;
    END
  END la1_data_out[3]
  PIN la1_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.580 4.000 145.780 ;
    END
  END la1_data_out[4]
  PIN la1_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.660 4.000 149.860 ;
    END
  END la1_data_out[5]
  PIN la1_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.740 4.000 153.940 ;
    END
  END la1_data_out[6]
  PIN la1_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.820 4.000 158.020 ;
    END
  END la1_data_out[7]
  PIN la1_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.900 4.000 162.100 ;
    END
  END la1_data_out[8]
  PIN la1_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.980 4.000 166.180 ;
    END
  END la1_data_out[9]
  PIN la1_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 1.100 300.000 2.300 ;
    END
  END la1_oenb[0]
  PIN la1_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 38.500 300.000 39.700 ;
    END
  END la1_oenb[10]
  PIN la1_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 41.900 300.000 43.100 ;
    END
  END la1_oenb[11]
  PIN la1_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 45.980 300.000 47.180 ;
    END
  END la1_oenb[12]
  PIN la1_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 49.380 300.000 50.580 ;
    END
  END la1_oenb[13]
  PIN la1_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 53.460 300.000 54.660 ;
    END
  END la1_oenb[14]
  PIN la1_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 56.860 300.000 58.060 ;
    END
  END la1_oenb[15]
  PIN la1_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 60.940 300.000 62.140 ;
    END
  END la1_oenb[16]
  PIN la1_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 64.340 300.000 65.540 ;
    END
  END la1_oenb[17]
  PIN la1_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 68.420 300.000 69.620 ;
    END
  END la1_oenb[18]
  PIN la1_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 71.820 300.000 73.020 ;
    END
  END la1_oenb[19]
  PIN la1_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 4.500 300.000 5.700 ;
    END
  END la1_oenb[1]
  PIN la1_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 75.900 300.000 77.100 ;
    END
  END la1_oenb[20]
  PIN la1_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 79.300 300.000 80.500 ;
    END
  END la1_oenb[21]
  PIN la1_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 83.380 300.000 84.580 ;
    END
  END la1_oenb[22]
  PIN la1_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 86.780 300.000 87.980 ;
    END
  END la1_oenb[23]
  PIN la1_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 90.860 300.000 92.060 ;
    END
  END la1_oenb[24]
  PIN la1_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 94.260 300.000 95.460 ;
    END
  END la1_oenb[25]
  PIN la1_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 98.340 300.000 99.540 ;
    END
  END la1_oenb[26]
  PIN la1_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 101.740 300.000 102.940 ;
    END
  END la1_oenb[27]
  PIN la1_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 105.820 300.000 107.020 ;
    END
  END la1_oenb[28]
  PIN la1_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 109.220 300.000 110.420 ;
    END
  END la1_oenb[29]
  PIN la1_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 8.580 300.000 9.780 ;
    END
  END la1_oenb[2]
  PIN la1_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 113.300 300.000 114.500 ;
    END
  END la1_oenb[30]
  PIN la1_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 116.700 300.000 117.900 ;
    END
  END la1_oenb[31]
  PIN la1_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 11.980 300.000 13.180 ;
    END
  END la1_oenb[3]
  PIN la1_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 16.060 300.000 17.260 ;
    END
  END la1_oenb[4]
  PIN la1_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 19.460 300.000 20.660 ;
    END
  END la1_oenb[5]
  PIN la1_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 23.540 300.000 24.740 ;
    END
  END la1_oenb[6]
  PIN la1_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 26.940 300.000 28.140 ;
    END
  END la1_oenb[7]
  PIN la1_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 31.020 300.000 32.220 ;
    END
  END la1_oenb[8]
  PIN la1_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 34.420 300.000 35.620 ;
    END
  END la1_oenb[9]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 2.480 22.640 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 2.480 176.240 288.560 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 2.480 99.440 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 2.480 253.040 288.560 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.610 296.000 10.170 300.000 ;
    END
  END wb_clk_i
  OBS
      LAYER li1 ;
        RECT 5.520 2.635 294.400 288.405 ;
      LAYER met1 ;
        RECT 3.290 2.480 296.630 289.980 ;
      LAYER met2 ;
        RECT 4.010 295.720 9.330 297.685 ;
        RECT 10.450 295.720 15.770 297.685 ;
        RECT 16.890 295.720 22.210 297.685 ;
        RECT 23.330 295.720 28.650 297.685 ;
        RECT 29.770 295.720 35.090 297.685 ;
        RECT 36.210 295.720 41.990 297.685 ;
        RECT 43.110 295.720 48.430 297.685 ;
        RECT 49.550 295.720 54.870 297.685 ;
        RECT 55.990 295.720 61.310 297.685 ;
        RECT 62.430 295.720 67.750 297.685 ;
        RECT 68.870 295.720 74.190 297.685 ;
        RECT 75.310 295.720 81.090 297.685 ;
        RECT 82.210 295.720 87.530 297.685 ;
        RECT 88.650 295.720 93.970 297.685 ;
        RECT 95.090 295.720 100.410 297.685 ;
        RECT 101.530 295.720 106.850 297.685 ;
        RECT 107.970 295.720 113.290 297.685 ;
        RECT 114.410 295.720 120.190 297.685 ;
        RECT 121.310 295.720 126.630 297.685 ;
        RECT 127.750 295.720 133.070 297.685 ;
        RECT 134.190 295.720 139.510 297.685 ;
        RECT 140.630 295.720 145.950 297.685 ;
        RECT 147.070 295.720 152.850 297.685 ;
        RECT 153.970 295.720 159.290 297.685 ;
        RECT 160.410 295.720 165.730 297.685 ;
        RECT 166.850 295.720 172.170 297.685 ;
        RECT 173.290 295.720 178.610 297.685 ;
        RECT 179.730 295.720 185.050 297.685 ;
        RECT 186.170 295.720 191.950 297.685 ;
        RECT 193.070 295.720 198.390 297.685 ;
        RECT 199.510 295.720 204.830 297.685 ;
        RECT 205.950 295.720 211.270 297.685 ;
        RECT 212.390 295.720 217.710 297.685 ;
        RECT 218.830 295.720 224.150 297.685 ;
        RECT 225.270 295.720 231.050 297.685 ;
        RECT 232.170 295.720 237.490 297.685 ;
        RECT 238.610 295.720 243.930 297.685 ;
        RECT 245.050 295.720 250.370 297.685 ;
        RECT 251.490 295.720 256.810 297.685 ;
        RECT 257.930 295.720 263.250 297.685 ;
        RECT 264.370 295.720 270.150 297.685 ;
        RECT 271.270 295.720 276.590 297.685 ;
        RECT 277.710 295.720 283.030 297.685 ;
        RECT 284.150 295.720 289.470 297.685 ;
        RECT 290.590 295.720 295.910 297.685 ;
        RECT 3.320 4.280 296.600 295.720 ;
        RECT 3.320 2.480 13.010 4.280 ;
        RECT 14.130 2.480 40.150 4.280 ;
        RECT 41.270 2.480 67.290 4.280 ;
        RECT 68.410 2.480 94.430 4.280 ;
        RECT 95.550 2.480 122.030 4.280 ;
        RECT 123.150 2.480 149.170 4.280 ;
        RECT 150.290 2.480 176.310 4.280 ;
        RECT 177.430 2.480 203.450 4.280 ;
        RECT 204.570 2.480 231.050 4.280 ;
        RECT 232.170 2.480 258.190 4.280 ;
        RECT 259.310 2.480 285.330 4.280 ;
        RECT 286.450 2.480 296.600 4.280 ;
      LAYER met3 ;
        RECT 4.400 296.500 295.600 297.665 ;
        RECT 4.000 294.420 296.000 296.500 ;
        RECT 4.400 292.420 295.600 294.420 ;
        RECT 4.000 291.020 296.000 292.420 ;
        RECT 4.000 290.340 295.600 291.020 ;
        RECT 4.400 289.020 295.600 290.340 ;
        RECT 4.400 288.340 296.000 289.020 ;
        RECT 4.000 286.940 296.000 288.340 ;
        RECT 4.000 286.260 295.600 286.940 ;
        RECT 4.400 284.940 295.600 286.260 ;
        RECT 4.400 284.260 296.000 284.940 ;
        RECT 4.000 283.540 296.000 284.260 ;
        RECT 4.000 282.180 295.600 283.540 ;
        RECT 4.400 281.540 295.600 282.180 ;
        RECT 4.400 280.180 296.000 281.540 ;
        RECT 4.000 279.460 296.000 280.180 ;
        RECT 4.000 278.100 295.600 279.460 ;
        RECT 4.400 277.460 295.600 278.100 ;
        RECT 4.400 276.100 296.000 277.460 ;
        RECT 4.000 276.060 296.000 276.100 ;
        RECT 4.000 274.060 295.600 276.060 ;
        RECT 4.000 274.020 296.000 274.060 ;
        RECT 4.400 272.020 296.000 274.020 ;
        RECT 4.000 271.980 296.000 272.020 ;
        RECT 4.000 269.980 295.600 271.980 ;
        RECT 4.000 269.940 296.000 269.980 ;
        RECT 4.400 268.580 296.000 269.940 ;
        RECT 4.400 267.940 295.600 268.580 ;
        RECT 4.000 266.580 295.600 267.940 ;
        RECT 4.000 266.540 296.000 266.580 ;
        RECT 4.400 264.540 296.000 266.540 ;
        RECT 4.000 264.500 296.000 264.540 ;
        RECT 4.000 262.500 295.600 264.500 ;
        RECT 4.000 262.460 296.000 262.500 ;
        RECT 4.400 261.100 296.000 262.460 ;
        RECT 4.400 260.460 295.600 261.100 ;
        RECT 4.000 259.100 295.600 260.460 ;
        RECT 4.000 258.380 296.000 259.100 ;
        RECT 4.400 257.020 296.000 258.380 ;
        RECT 4.400 256.380 295.600 257.020 ;
        RECT 4.000 255.020 295.600 256.380 ;
        RECT 4.000 254.300 296.000 255.020 ;
        RECT 4.400 253.620 296.000 254.300 ;
        RECT 4.400 252.300 295.600 253.620 ;
        RECT 4.000 251.620 295.600 252.300 ;
        RECT 4.000 250.220 296.000 251.620 ;
        RECT 4.400 249.540 296.000 250.220 ;
        RECT 4.400 248.220 295.600 249.540 ;
        RECT 4.000 247.540 295.600 248.220 ;
        RECT 4.000 246.140 296.000 247.540 ;
        RECT 4.400 244.140 295.600 246.140 ;
        RECT 4.000 242.060 296.000 244.140 ;
        RECT 4.400 240.060 295.600 242.060 ;
        RECT 4.000 238.660 296.000 240.060 ;
        RECT 4.000 237.980 295.600 238.660 ;
        RECT 4.400 236.660 295.600 237.980 ;
        RECT 4.400 235.980 296.000 236.660 ;
        RECT 4.000 234.580 296.000 235.980 ;
        RECT 4.400 232.580 295.600 234.580 ;
        RECT 4.000 231.180 296.000 232.580 ;
        RECT 4.000 230.500 295.600 231.180 ;
        RECT 4.400 229.180 295.600 230.500 ;
        RECT 4.400 228.500 296.000 229.180 ;
        RECT 4.000 227.100 296.000 228.500 ;
        RECT 4.000 226.420 295.600 227.100 ;
        RECT 4.400 225.100 295.600 226.420 ;
        RECT 4.400 224.420 296.000 225.100 ;
        RECT 4.000 223.700 296.000 224.420 ;
        RECT 4.000 222.340 295.600 223.700 ;
        RECT 4.400 221.700 295.600 222.340 ;
        RECT 4.400 220.340 296.000 221.700 ;
        RECT 4.000 219.620 296.000 220.340 ;
        RECT 4.000 218.260 295.600 219.620 ;
        RECT 4.400 217.620 295.600 218.260 ;
        RECT 4.400 216.260 296.000 217.620 ;
        RECT 4.000 216.220 296.000 216.260 ;
        RECT 4.000 214.220 295.600 216.220 ;
        RECT 4.000 214.180 296.000 214.220 ;
        RECT 4.400 212.180 296.000 214.180 ;
        RECT 4.000 212.140 296.000 212.180 ;
        RECT 4.000 210.140 295.600 212.140 ;
        RECT 4.000 210.100 296.000 210.140 ;
        RECT 4.400 208.740 296.000 210.100 ;
        RECT 4.400 208.100 295.600 208.740 ;
        RECT 4.000 206.740 295.600 208.100 ;
        RECT 4.000 206.020 296.000 206.740 ;
        RECT 4.400 204.660 296.000 206.020 ;
        RECT 4.400 204.020 295.600 204.660 ;
        RECT 4.000 202.660 295.600 204.020 ;
        RECT 4.000 202.620 296.000 202.660 ;
        RECT 4.400 201.260 296.000 202.620 ;
        RECT 4.400 200.620 295.600 201.260 ;
        RECT 4.000 199.260 295.600 200.620 ;
        RECT 4.000 198.540 296.000 199.260 ;
        RECT 4.400 197.180 296.000 198.540 ;
        RECT 4.400 196.540 295.600 197.180 ;
        RECT 4.000 195.180 295.600 196.540 ;
        RECT 4.000 194.460 296.000 195.180 ;
        RECT 4.400 193.780 296.000 194.460 ;
        RECT 4.400 192.460 295.600 193.780 ;
        RECT 4.000 191.780 295.600 192.460 ;
        RECT 4.000 190.380 296.000 191.780 ;
        RECT 4.400 189.700 296.000 190.380 ;
        RECT 4.400 188.380 295.600 189.700 ;
        RECT 4.000 187.700 295.600 188.380 ;
        RECT 4.000 186.300 296.000 187.700 ;
        RECT 4.400 184.300 295.600 186.300 ;
        RECT 4.000 182.220 296.000 184.300 ;
        RECT 4.400 180.220 295.600 182.220 ;
        RECT 4.000 178.820 296.000 180.220 ;
        RECT 4.000 178.140 295.600 178.820 ;
        RECT 4.400 176.820 295.600 178.140 ;
        RECT 4.400 176.140 296.000 176.820 ;
        RECT 4.000 174.740 296.000 176.140 ;
        RECT 4.000 174.060 295.600 174.740 ;
        RECT 4.400 172.740 295.600 174.060 ;
        RECT 4.400 172.060 296.000 172.740 ;
        RECT 4.000 171.340 296.000 172.060 ;
        RECT 4.000 169.980 295.600 171.340 ;
        RECT 4.400 169.340 295.600 169.980 ;
        RECT 4.400 167.980 296.000 169.340 ;
        RECT 4.000 167.260 296.000 167.980 ;
        RECT 4.000 166.580 295.600 167.260 ;
        RECT 4.400 165.260 295.600 166.580 ;
        RECT 4.400 164.580 296.000 165.260 ;
        RECT 4.000 163.860 296.000 164.580 ;
        RECT 4.000 162.500 295.600 163.860 ;
        RECT 4.400 161.860 295.600 162.500 ;
        RECT 4.400 160.500 296.000 161.860 ;
        RECT 4.000 159.780 296.000 160.500 ;
        RECT 4.000 158.420 295.600 159.780 ;
        RECT 4.400 157.780 295.600 158.420 ;
        RECT 4.400 156.420 296.000 157.780 ;
        RECT 4.000 156.380 296.000 156.420 ;
        RECT 4.000 154.380 295.600 156.380 ;
        RECT 4.000 154.340 296.000 154.380 ;
        RECT 4.400 152.340 296.000 154.340 ;
        RECT 4.000 152.300 296.000 152.340 ;
        RECT 4.000 150.300 295.600 152.300 ;
        RECT 4.000 150.260 296.000 150.300 ;
        RECT 4.400 148.260 296.000 150.260 ;
        RECT 4.000 148.220 296.000 148.260 ;
        RECT 4.000 146.220 295.600 148.220 ;
        RECT 4.000 146.180 296.000 146.220 ;
        RECT 4.400 144.820 296.000 146.180 ;
        RECT 4.400 144.180 295.600 144.820 ;
        RECT 4.000 142.820 295.600 144.180 ;
        RECT 4.000 142.100 296.000 142.820 ;
        RECT 4.400 140.740 296.000 142.100 ;
        RECT 4.400 140.100 295.600 140.740 ;
        RECT 4.000 138.740 295.600 140.100 ;
        RECT 4.000 138.020 296.000 138.740 ;
        RECT 4.400 137.340 296.000 138.020 ;
        RECT 4.400 136.020 295.600 137.340 ;
        RECT 4.000 135.340 295.600 136.020 ;
        RECT 4.000 134.620 296.000 135.340 ;
        RECT 4.400 133.260 296.000 134.620 ;
        RECT 4.400 132.620 295.600 133.260 ;
        RECT 4.000 131.260 295.600 132.620 ;
        RECT 4.000 130.540 296.000 131.260 ;
        RECT 4.400 129.860 296.000 130.540 ;
        RECT 4.400 128.540 295.600 129.860 ;
        RECT 4.000 127.860 295.600 128.540 ;
        RECT 4.000 126.460 296.000 127.860 ;
        RECT 4.400 125.780 296.000 126.460 ;
        RECT 4.400 124.460 295.600 125.780 ;
        RECT 4.000 123.780 295.600 124.460 ;
        RECT 4.000 122.380 296.000 123.780 ;
        RECT 4.400 120.380 295.600 122.380 ;
        RECT 4.000 118.300 296.000 120.380 ;
        RECT 4.400 116.300 295.600 118.300 ;
        RECT 4.000 114.900 296.000 116.300 ;
        RECT 4.000 114.220 295.600 114.900 ;
        RECT 4.400 112.900 295.600 114.220 ;
        RECT 4.400 112.220 296.000 112.900 ;
        RECT 4.000 110.820 296.000 112.220 ;
        RECT 4.000 110.140 295.600 110.820 ;
        RECT 4.400 108.820 295.600 110.140 ;
        RECT 4.400 108.140 296.000 108.820 ;
        RECT 4.000 107.420 296.000 108.140 ;
        RECT 4.000 106.060 295.600 107.420 ;
        RECT 4.400 105.420 295.600 106.060 ;
        RECT 4.400 104.060 296.000 105.420 ;
        RECT 4.000 103.340 296.000 104.060 ;
        RECT 4.000 102.660 295.600 103.340 ;
        RECT 4.400 101.340 295.600 102.660 ;
        RECT 4.400 100.660 296.000 101.340 ;
        RECT 4.000 99.940 296.000 100.660 ;
        RECT 4.000 98.580 295.600 99.940 ;
        RECT 4.400 97.940 295.600 98.580 ;
        RECT 4.400 96.580 296.000 97.940 ;
        RECT 4.000 95.860 296.000 96.580 ;
        RECT 4.000 94.500 295.600 95.860 ;
        RECT 4.400 93.860 295.600 94.500 ;
        RECT 4.400 92.500 296.000 93.860 ;
        RECT 4.000 92.460 296.000 92.500 ;
        RECT 4.000 90.460 295.600 92.460 ;
        RECT 4.000 90.420 296.000 90.460 ;
        RECT 4.400 88.420 296.000 90.420 ;
        RECT 4.000 88.380 296.000 88.420 ;
        RECT 4.000 86.380 295.600 88.380 ;
        RECT 4.000 86.340 296.000 86.380 ;
        RECT 4.400 84.980 296.000 86.340 ;
        RECT 4.400 84.340 295.600 84.980 ;
        RECT 4.000 82.980 295.600 84.340 ;
        RECT 4.000 82.260 296.000 82.980 ;
        RECT 4.400 80.900 296.000 82.260 ;
        RECT 4.400 80.260 295.600 80.900 ;
        RECT 4.000 78.900 295.600 80.260 ;
        RECT 4.000 78.180 296.000 78.900 ;
        RECT 4.400 77.500 296.000 78.180 ;
        RECT 4.400 76.180 295.600 77.500 ;
        RECT 4.000 75.500 295.600 76.180 ;
        RECT 4.000 74.100 296.000 75.500 ;
        RECT 4.400 73.420 296.000 74.100 ;
        RECT 4.400 72.100 295.600 73.420 ;
        RECT 4.000 71.420 295.600 72.100 ;
        RECT 4.000 70.020 296.000 71.420 ;
        RECT 4.400 68.020 295.600 70.020 ;
        RECT 4.000 66.620 296.000 68.020 ;
        RECT 4.400 65.940 296.000 66.620 ;
        RECT 4.400 64.620 295.600 65.940 ;
        RECT 4.000 63.940 295.600 64.620 ;
        RECT 4.000 62.540 296.000 63.940 ;
        RECT 4.400 60.540 295.600 62.540 ;
        RECT 4.000 58.460 296.000 60.540 ;
        RECT 4.400 56.460 295.600 58.460 ;
        RECT 4.000 55.060 296.000 56.460 ;
        RECT 4.000 54.380 295.600 55.060 ;
        RECT 4.400 53.060 295.600 54.380 ;
        RECT 4.400 52.380 296.000 53.060 ;
        RECT 4.000 50.980 296.000 52.380 ;
        RECT 4.000 50.300 295.600 50.980 ;
        RECT 4.400 48.980 295.600 50.300 ;
        RECT 4.400 48.300 296.000 48.980 ;
        RECT 4.000 47.580 296.000 48.300 ;
        RECT 4.000 46.220 295.600 47.580 ;
        RECT 4.400 45.580 295.600 46.220 ;
        RECT 4.400 44.220 296.000 45.580 ;
        RECT 4.000 43.500 296.000 44.220 ;
        RECT 4.000 42.140 295.600 43.500 ;
        RECT 4.400 41.500 295.600 42.140 ;
        RECT 4.400 40.140 296.000 41.500 ;
        RECT 4.000 40.100 296.000 40.140 ;
        RECT 4.000 38.100 295.600 40.100 ;
        RECT 4.000 38.060 296.000 38.100 ;
        RECT 4.400 36.060 296.000 38.060 ;
        RECT 4.000 36.020 296.000 36.060 ;
        RECT 4.000 34.660 295.600 36.020 ;
        RECT 4.400 34.020 295.600 34.660 ;
        RECT 4.400 32.660 296.000 34.020 ;
        RECT 4.000 32.620 296.000 32.660 ;
        RECT 4.000 30.620 295.600 32.620 ;
        RECT 4.000 30.580 296.000 30.620 ;
        RECT 4.400 28.580 296.000 30.580 ;
        RECT 4.000 28.540 296.000 28.580 ;
        RECT 4.000 26.540 295.600 28.540 ;
        RECT 4.000 26.500 296.000 26.540 ;
        RECT 4.400 25.140 296.000 26.500 ;
        RECT 4.400 24.500 295.600 25.140 ;
        RECT 4.000 23.140 295.600 24.500 ;
        RECT 4.000 22.420 296.000 23.140 ;
        RECT 4.400 21.060 296.000 22.420 ;
        RECT 4.400 20.420 295.600 21.060 ;
        RECT 4.000 19.060 295.600 20.420 ;
        RECT 4.000 18.340 296.000 19.060 ;
        RECT 4.400 17.660 296.000 18.340 ;
        RECT 4.400 16.340 295.600 17.660 ;
        RECT 4.000 15.660 295.600 16.340 ;
        RECT 4.000 14.260 296.000 15.660 ;
        RECT 4.400 13.580 296.000 14.260 ;
        RECT 4.400 12.260 295.600 13.580 ;
        RECT 4.000 11.580 295.600 12.260 ;
        RECT 4.000 10.180 296.000 11.580 ;
        RECT 4.400 8.180 295.600 10.180 ;
        RECT 4.000 6.100 296.000 8.180 ;
        RECT 4.400 4.100 295.600 6.100 ;
        RECT 4.000 2.700 296.000 4.100 ;
        RECT 4.400 2.555 295.600 2.700 ;
      LAYER met4 ;
        RECT 23.295 6.975 97.440 272.505 ;
        RECT 99.840 6.975 174.240 272.505 ;
        RECT 176.640 6.975 249.945 272.505 ;
  END
END wrapped_vgademo_on_fpga
END LIBRARY

