VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_vgademo_on_fpga
  CLASS BLOCK ;
  FOREIGN wrapped_vgademo_on_fpga ;
  ORIGIN 0.000 0.000 ;
  SIZE 300.000 BY 280.000 ;
  PIN active
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.710 276.000 3.270 280.000 ;
    END
  END active
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.750 276.000 14.310 280.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.950 276.000 69.510 280.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.470 276.000 75.030 280.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.450 276.000 81.010 280.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.970 276.000 86.530 280.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.490 276.000 92.050 280.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.010 276.000 97.570 280.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.530 276.000 103.090 280.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.050 276.000 108.610 280.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.570 276.000 114.130 280.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.090 276.000 119.650 280.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.270 276.000 19.830 280.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.610 276.000 125.170 280.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.130 276.000 130.690 280.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.650 276.000 136.210 280.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.170 276.000 141.730 280.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.690 276.000 147.250 280.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.670 276.000 153.230 280.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.190 276.000 158.750 280.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.710 276.000 164.270 280.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.230 276.000 169.790 280.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.750 276.000 175.310 280.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.790 276.000 25.350 280.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.270 276.000 180.830 280.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.790 276.000 186.350 280.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.310 276.000 191.870 280.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.830 276.000 197.390 280.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.350 276.000 202.910 280.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.870 276.000 208.430 280.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.390 276.000 213.950 280.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.910 276.000 219.470 280.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.310 276.000 30.870 280.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.830 276.000 36.390 280.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.350 276.000 41.910 280.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.870 276.000 47.430 280.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.390 276.000 52.950 280.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.910 276.000 58.470 280.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.430 276.000 63.990 280.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 111.260 300.000 112.460 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 145.940 300.000 147.140 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 149.340 300.000 150.540 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 152.740 300.000 153.940 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 156.140 300.000 157.340 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 159.540 300.000 160.740 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 163.620 300.000 164.820 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 167.020 300.000 168.220 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 170.420 300.000 171.620 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 173.820 300.000 175.020 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 177.220 300.000 178.420 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 114.660 300.000 115.860 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 180.620 300.000 181.820 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 184.020 300.000 185.220 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 187.420 300.000 188.620 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 190.820 300.000 192.020 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 194.220 300.000 195.420 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 197.620 300.000 198.820 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 201.700 300.000 202.900 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 205.100 300.000 206.300 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 208.500 300.000 209.700 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 211.900 300.000 213.100 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 118.060 300.000 119.260 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 215.300 300.000 216.500 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 218.700 300.000 219.900 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 222.100 300.000 223.300 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 225.500 300.000 226.700 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 228.900 300.000 230.100 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 232.300 300.000 233.500 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 235.700 300.000 236.900 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 239.100 300.000 240.300 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 122.140 300.000 123.340 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 125.540 300.000 126.740 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 128.940 300.000 130.140 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 132.340 300.000 133.540 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 135.740 300.000 136.940 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 139.140 300.000 140.340 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 142.540 300.000 143.740 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 243.180 300.000 244.380 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 253.380 300.000 254.580 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 256.780 300.000 257.980 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.610 0.000 56.170 4.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.490 276.000 253.050 280.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.330 0.000 93.890 4.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.590 0.000 131.150 4.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.310 0.000 168.870 4.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.010 276.000 258.570 280.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 260.180 300.000 261.380 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 263.580 300.000 264.780 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 260.860 4.000 262.060 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.530 276.000 264.090 280.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 264.940 4.000 266.140 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 266.980 300.000 268.180 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.050 276.000 269.610 280.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 270.380 300.000 271.580 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 273.780 300.000 274.980 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 269.020 4.000 270.220 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.570 276.000 275.130 280.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.090 276.000 280.650 280.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.610 276.000 286.170 280.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.430 276.000 224.990 280.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.130 276.000 291.690 280.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.570 0.000 206.130 4.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 277.180 300.000 278.380 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.290 0.000 243.850 4.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.550 0.000 281.110 4.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 273.100 4.000 274.300 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.650 276.000 297.210 280.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 277.180 4.000 278.380 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.410 276.000 230.970 280.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.930 276.000 236.490 280.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.350 0.000 18.910 4.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.450 276.000 242.010 280.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 246.580 300.000 247.780 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 249.980 300.000 251.180 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.970 276.000 247.530 280.000 ;
    END
  END io_out[9]
  PIN la1_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1.100 4.000 2.300 ;
    END
  END la1_data_in[0]
  PIN la1_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 41.220 4.000 42.420 ;
    END
  END la1_data_in[10]
  PIN la1_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.300 4.000 46.500 ;
    END
  END la1_data_in[11]
  PIN la1_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.380 4.000 50.580 ;
    END
  END la1_data_in[12]
  PIN la1_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.460 4.000 54.660 ;
    END
  END la1_data_in[13]
  PIN la1_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.540 4.000 58.740 ;
    END
  END la1_data_in[14]
  PIN la1_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.620 4.000 62.820 ;
    END
  END la1_data_in[15]
  PIN la1_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.700 4.000 66.900 ;
    END
  END la1_data_in[16]
  PIN la1_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.780 4.000 70.980 ;
    END
  END la1_data_in[17]
  PIN la1_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.860 4.000 75.060 ;
    END
  END la1_data_in[18]
  PIN la1_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.940 4.000 79.140 ;
    END
  END la1_data_in[19]
  PIN la1_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.500 4.000 5.700 ;
    END
  END la1_data_in[1]
  PIN la1_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 82.020 4.000 83.220 ;
    END
  END la1_data_in[20]
  PIN la1_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 86.100 4.000 87.300 ;
    END
  END la1_data_in[21]
  PIN la1_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 90.180 4.000 91.380 ;
    END
  END la1_data_in[22]
  PIN la1_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 94.260 4.000 95.460 ;
    END
  END la1_data_in[23]
  PIN la1_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.340 4.000 99.540 ;
    END
  END la1_data_in[24]
  PIN la1_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.420 4.000 103.620 ;
    END
  END la1_data_in[25]
  PIN la1_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.500 4.000 107.700 ;
    END
  END la1_data_in[26]
  PIN la1_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.580 4.000 111.780 ;
    END
  END la1_data_in[27]
  PIN la1_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.660 4.000 115.860 ;
    END
  END la1_data_in[28]
  PIN la1_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.740 4.000 119.940 ;
    END
  END la1_data_in[29]
  PIN la1_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.580 4.000 9.780 ;
    END
  END la1_data_in[2]
  PIN la1_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.820 4.000 124.020 ;
    END
  END la1_data_in[30]
  PIN la1_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.900 4.000 128.100 ;
    END
  END la1_data_in[31]
  PIN la1_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.660 4.000 13.860 ;
    END
  END la1_data_in[3]
  PIN la1_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.740 4.000 17.940 ;
    END
  END la1_data_in[4]
  PIN la1_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.820 4.000 22.020 ;
    END
  END la1_data_in[5]
  PIN la1_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.900 4.000 26.100 ;
    END
  END la1_data_in[6]
  PIN la1_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.980 4.000 30.180 ;
    END
  END la1_data_in[7]
  PIN la1_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.060 4.000 34.260 ;
    END
  END la1_data_in[8]
  PIN la1_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.140 4.000 38.340 ;
    END
  END la1_data_in[9]
  PIN la1_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.980 4.000 132.180 ;
    END
  END la1_data_out[0]
  PIN la1_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 171.100 4.000 172.300 ;
    END
  END la1_data_out[10]
  PIN la1_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.180 4.000 176.380 ;
    END
  END la1_data_out[11]
  PIN la1_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.260 4.000 180.460 ;
    END
  END la1_data_out[12]
  PIN la1_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.340 4.000 184.540 ;
    END
  END la1_data_out[13]
  PIN la1_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.420 4.000 188.620 ;
    END
  END la1_data_out[14]
  PIN la1_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.500 4.000 192.700 ;
    END
  END la1_data_out[15]
  PIN la1_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.580 4.000 196.780 ;
    END
  END la1_data_out[16]
  PIN la1_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.660 4.000 200.860 ;
    END
  END la1_data_out[17]
  PIN la1_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 203.740 4.000 204.940 ;
    END
  END la1_data_out[18]
  PIN la1_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.820 4.000 209.020 ;
    END
  END la1_data_out[19]
  PIN la1_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 135.060 4.000 136.260 ;
    END
  END la1_data_out[1]
  PIN la1_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 211.900 4.000 213.100 ;
    END
  END la1_data_out[20]
  PIN la1_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 215.980 4.000 217.180 ;
    END
  END la1_data_out[21]
  PIN la1_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 220.060 4.000 221.260 ;
    END
  END la1_data_out[22]
  PIN la1_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.140 4.000 225.340 ;
    END
  END la1_data_out[23]
  PIN la1_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 228.220 4.000 229.420 ;
    END
  END la1_data_out[24]
  PIN la1_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 232.300 4.000 233.500 ;
    END
  END la1_data_out[25]
  PIN la1_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.380 4.000 237.580 ;
    END
  END la1_data_out[26]
  PIN la1_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.460 4.000 241.660 ;
    END
  END la1_data_out[27]
  PIN la1_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.540 4.000 245.740 ;
    END
  END la1_data_out[28]
  PIN la1_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.620 4.000 249.820 ;
    END
  END la1_data_out[29]
  PIN la1_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.140 4.000 140.340 ;
    END
  END la1_data_out[2]
  PIN la1_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 252.700 4.000 253.900 ;
    END
  END la1_data_out[30]
  PIN la1_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 256.780 4.000 257.980 ;
    END
  END la1_data_out[31]
  PIN la1_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.540 4.000 143.740 ;
    END
  END la1_data_out[3]
  PIN la1_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.620 4.000 147.820 ;
    END
  END la1_data_out[4]
  PIN la1_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 150.700 4.000 151.900 ;
    END
  END la1_data_out[5]
  PIN la1_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 154.780 4.000 155.980 ;
    END
  END la1_data_out[6]
  PIN la1_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 158.860 4.000 160.060 ;
    END
  END la1_data_out[7]
  PIN la1_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 162.940 4.000 164.140 ;
    END
  END la1_data_out[8]
  PIN la1_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 167.020 4.000 168.220 ;
    END
  END la1_data_out[9]
  PIN la1_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 1.100 300.000 2.300 ;
    END
  END la1_oenb[0]
  PIN la1_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 35.100 300.000 36.300 ;
    END
  END la1_oenb[10]
  PIN la1_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 38.500 300.000 39.700 ;
    END
  END la1_oenb[11]
  PIN la1_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 42.580 300.000 43.780 ;
    END
  END la1_oenb[12]
  PIN la1_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 45.980 300.000 47.180 ;
    END
  END la1_oenb[13]
  PIN la1_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 49.380 300.000 50.580 ;
    END
  END la1_oenb[14]
  PIN la1_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 52.780 300.000 53.980 ;
    END
  END la1_oenb[15]
  PIN la1_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 56.180 300.000 57.380 ;
    END
  END la1_oenb[16]
  PIN la1_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 59.580 300.000 60.780 ;
    END
  END la1_oenb[17]
  PIN la1_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 62.980 300.000 64.180 ;
    END
  END la1_oenb[18]
  PIN la1_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 66.380 300.000 67.580 ;
    END
  END la1_oenb[19]
  PIN la1_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 4.500 300.000 5.700 ;
    END
  END la1_oenb[1]
  PIN la1_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 69.780 300.000 70.980 ;
    END
  END la1_oenb[20]
  PIN la1_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 73.180 300.000 74.380 ;
    END
  END la1_oenb[21]
  PIN la1_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 76.580 300.000 77.780 ;
    END
  END la1_oenb[22]
  PIN la1_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 79.980 300.000 81.180 ;
    END
  END la1_oenb[23]
  PIN la1_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 84.060 300.000 85.260 ;
    END
  END la1_oenb[24]
  PIN la1_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 87.460 300.000 88.660 ;
    END
  END la1_oenb[25]
  PIN la1_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 90.860 300.000 92.060 ;
    END
  END la1_oenb[26]
  PIN la1_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 94.260 300.000 95.460 ;
    END
  END la1_oenb[27]
  PIN la1_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 97.660 300.000 98.860 ;
    END
  END la1_oenb[28]
  PIN la1_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 101.060 300.000 102.260 ;
    END
  END la1_oenb[29]
  PIN la1_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 7.900 300.000 9.100 ;
    END
  END la1_oenb[2]
  PIN la1_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 104.460 300.000 105.660 ;
    END
  END la1_oenb[30]
  PIN la1_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 107.860 300.000 109.060 ;
    END
  END la1_oenb[31]
  PIN la1_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 11.300 300.000 12.500 ;
    END
  END la1_oenb[3]
  PIN la1_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 14.700 300.000 15.900 ;
    END
  END la1_oenb[4]
  PIN la1_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 18.100 300.000 19.300 ;
    END
  END la1_oenb[5]
  PIN la1_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 21.500 300.000 22.700 ;
    END
  END la1_oenb[6]
  PIN la1_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 24.900 300.000 26.100 ;
    END
  END la1_oenb[7]
  PIN la1_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 28.300 300.000 29.500 ;
    END
  END la1_oenb[8]
  PIN la1_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 31.700 300.000 32.900 ;
    END
  END la1_oenb[9]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 2.480 22.640 266.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 2.480 176.240 266.800 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 2.480 99.440 266.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 2.480 253.040 266.800 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.230 276.000 8.790 280.000 ;
    END
  END wb_clk_i
  OBS
      LAYER li1 ;
        RECT 5.520 2.635 294.400 266.645 ;
      LAYER met1 ;
        RECT 2.830 1.400 297.090 269.240 ;
      LAYER met2 ;
        RECT 3.550 275.720 7.950 277.965 ;
        RECT 9.070 275.720 13.470 277.965 ;
        RECT 14.590 275.720 18.990 277.965 ;
        RECT 20.110 275.720 24.510 277.965 ;
        RECT 25.630 275.720 30.030 277.965 ;
        RECT 31.150 275.720 35.550 277.965 ;
        RECT 36.670 275.720 41.070 277.965 ;
        RECT 42.190 275.720 46.590 277.965 ;
        RECT 47.710 275.720 52.110 277.965 ;
        RECT 53.230 275.720 57.630 277.965 ;
        RECT 58.750 275.720 63.150 277.965 ;
        RECT 64.270 275.720 68.670 277.965 ;
        RECT 69.790 275.720 74.190 277.965 ;
        RECT 75.310 275.720 80.170 277.965 ;
        RECT 81.290 275.720 85.690 277.965 ;
        RECT 86.810 275.720 91.210 277.965 ;
        RECT 92.330 275.720 96.730 277.965 ;
        RECT 97.850 275.720 102.250 277.965 ;
        RECT 103.370 275.720 107.770 277.965 ;
        RECT 108.890 275.720 113.290 277.965 ;
        RECT 114.410 275.720 118.810 277.965 ;
        RECT 119.930 275.720 124.330 277.965 ;
        RECT 125.450 275.720 129.850 277.965 ;
        RECT 130.970 275.720 135.370 277.965 ;
        RECT 136.490 275.720 140.890 277.965 ;
        RECT 142.010 275.720 146.410 277.965 ;
        RECT 147.530 275.720 152.390 277.965 ;
        RECT 153.510 275.720 157.910 277.965 ;
        RECT 159.030 275.720 163.430 277.965 ;
        RECT 164.550 275.720 168.950 277.965 ;
        RECT 170.070 275.720 174.470 277.965 ;
        RECT 175.590 275.720 179.990 277.965 ;
        RECT 181.110 275.720 185.510 277.965 ;
        RECT 186.630 275.720 191.030 277.965 ;
        RECT 192.150 275.720 196.550 277.965 ;
        RECT 197.670 275.720 202.070 277.965 ;
        RECT 203.190 275.720 207.590 277.965 ;
        RECT 208.710 275.720 213.110 277.965 ;
        RECT 214.230 275.720 218.630 277.965 ;
        RECT 219.750 275.720 224.150 277.965 ;
        RECT 225.270 275.720 230.130 277.965 ;
        RECT 231.250 275.720 235.650 277.965 ;
        RECT 236.770 275.720 241.170 277.965 ;
        RECT 242.290 275.720 246.690 277.965 ;
        RECT 247.810 275.720 252.210 277.965 ;
        RECT 253.330 275.720 257.730 277.965 ;
        RECT 258.850 275.720 263.250 277.965 ;
        RECT 264.370 275.720 268.770 277.965 ;
        RECT 269.890 275.720 274.290 277.965 ;
        RECT 275.410 275.720 279.810 277.965 ;
        RECT 280.930 275.720 285.330 277.965 ;
        RECT 286.450 275.720 290.850 277.965 ;
        RECT 291.970 275.720 296.370 277.965 ;
        RECT 2.860 4.280 297.060 275.720 ;
        RECT 2.860 1.370 18.070 4.280 ;
        RECT 19.190 1.370 55.330 4.280 ;
        RECT 56.450 1.370 93.050 4.280 ;
        RECT 94.170 1.370 130.310 4.280 ;
        RECT 131.430 1.370 168.030 4.280 ;
        RECT 169.150 1.370 205.290 4.280 ;
        RECT 206.410 1.370 243.010 4.280 ;
        RECT 244.130 1.370 280.270 4.280 ;
        RECT 281.390 1.370 297.060 4.280 ;
      LAYER met3 ;
        RECT 4.400 276.780 295.600 277.945 ;
        RECT 4.000 275.380 296.000 276.780 ;
        RECT 4.000 274.700 295.600 275.380 ;
        RECT 4.400 273.380 295.600 274.700 ;
        RECT 4.400 272.700 296.000 273.380 ;
        RECT 4.000 271.980 296.000 272.700 ;
        RECT 4.000 270.620 295.600 271.980 ;
        RECT 4.400 269.980 295.600 270.620 ;
        RECT 4.400 268.620 296.000 269.980 ;
        RECT 4.000 268.580 296.000 268.620 ;
        RECT 4.000 266.580 295.600 268.580 ;
        RECT 4.000 266.540 296.000 266.580 ;
        RECT 4.400 265.180 296.000 266.540 ;
        RECT 4.400 264.540 295.600 265.180 ;
        RECT 4.000 263.180 295.600 264.540 ;
        RECT 4.000 262.460 296.000 263.180 ;
        RECT 4.400 261.780 296.000 262.460 ;
        RECT 4.400 260.460 295.600 261.780 ;
        RECT 4.000 259.780 295.600 260.460 ;
        RECT 4.000 258.380 296.000 259.780 ;
        RECT 4.400 256.380 295.600 258.380 ;
        RECT 4.000 254.980 296.000 256.380 ;
        RECT 4.000 254.300 295.600 254.980 ;
        RECT 4.400 252.980 295.600 254.300 ;
        RECT 4.400 252.300 296.000 252.980 ;
        RECT 4.000 251.580 296.000 252.300 ;
        RECT 4.000 250.220 295.600 251.580 ;
        RECT 4.400 249.580 295.600 250.220 ;
        RECT 4.400 248.220 296.000 249.580 ;
        RECT 4.000 248.180 296.000 248.220 ;
        RECT 4.000 246.180 295.600 248.180 ;
        RECT 4.000 246.140 296.000 246.180 ;
        RECT 4.400 244.780 296.000 246.140 ;
        RECT 4.400 244.140 295.600 244.780 ;
        RECT 4.000 242.780 295.600 244.140 ;
        RECT 4.000 242.060 296.000 242.780 ;
        RECT 4.400 240.700 296.000 242.060 ;
        RECT 4.400 240.060 295.600 240.700 ;
        RECT 4.000 238.700 295.600 240.060 ;
        RECT 4.000 237.980 296.000 238.700 ;
        RECT 4.400 237.300 296.000 237.980 ;
        RECT 4.400 235.980 295.600 237.300 ;
        RECT 4.000 235.300 295.600 235.980 ;
        RECT 4.000 233.900 296.000 235.300 ;
        RECT 4.400 231.900 295.600 233.900 ;
        RECT 4.000 230.500 296.000 231.900 ;
        RECT 4.000 229.820 295.600 230.500 ;
        RECT 4.400 228.500 295.600 229.820 ;
        RECT 4.400 227.820 296.000 228.500 ;
        RECT 4.000 227.100 296.000 227.820 ;
        RECT 4.000 225.740 295.600 227.100 ;
        RECT 4.400 225.100 295.600 225.740 ;
        RECT 4.400 223.740 296.000 225.100 ;
        RECT 4.000 223.700 296.000 223.740 ;
        RECT 4.000 221.700 295.600 223.700 ;
        RECT 4.000 221.660 296.000 221.700 ;
        RECT 4.400 220.300 296.000 221.660 ;
        RECT 4.400 219.660 295.600 220.300 ;
        RECT 4.000 218.300 295.600 219.660 ;
        RECT 4.000 217.580 296.000 218.300 ;
        RECT 4.400 216.900 296.000 217.580 ;
        RECT 4.400 215.580 295.600 216.900 ;
        RECT 4.000 214.900 295.600 215.580 ;
        RECT 4.000 213.500 296.000 214.900 ;
        RECT 4.400 211.500 295.600 213.500 ;
        RECT 4.000 210.100 296.000 211.500 ;
        RECT 4.000 209.420 295.600 210.100 ;
        RECT 4.400 208.100 295.600 209.420 ;
        RECT 4.400 207.420 296.000 208.100 ;
        RECT 4.000 206.700 296.000 207.420 ;
        RECT 4.000 205.340 295.600 206.700 ;
        RECT 4.400 204.700 295.600 205.340 ;
        RECT 4.400 203.340 296.000 204.700 ;
        RECT 4.000 203.300 296.000 203.340 ;
        RECT 4.000 201.300 295.600 203.300 ;
        RECT 4.000 201.260 296.000 201.300 ;
        RECT 4.400 199.260 296.000 201.260 ;
        RECT 4.000 199.220 296.000 199.260 ;
        RECT 4.000 197.220 295.600 199.220 ;
        RECT 4.000 197.180 296.000 197.220 ;
        RECT 4.400 195.820 296.000 197.180 ;
        RECT 4.400 195.180 295.600 195.820 ;
        RECT 4.000 193.820 295.600 195.180 ;
        RECT 4.000 193.100 296.000 193.820 ;
        RECT 4.400 192.420 296.000 193.100 ;
        RECT 4.400 191.100 295.600 192.420 ;
        RECT 4.000 190.420 295.600 191.100 ;
        RECT 4.000 189.020 296.000 190.420 ;
        RECT 4.400 187.020 295.600 189.020 ;
        RECT 4.000 185.620 296.000 187.020 ;
        RECT 4.000 184.940 295.600 185.620 ;
        RECT 4.400 183.620 295.600 184.940 ;
        RECT 4.400 182.940 296.000 183.620 ;
        RECT 4.000 182.220 296.000 182.940 ;
        RECT 4.000 180.860 295.600 182.220 ;
        RECT 4.400 180.220 295.600 180.860 ;
        RECT 4.400 178.860 296.000 180.220 ;
        RECT 4.000 178.820 296.000 178.860 ;
        RECT 4.000 176.820 295.600 178.820 ;
        RECT 4.000 176.780 296.000 176.820 ;
        RECT 4.400 175.420 296.000 176.780 ;
        RECT 4.400 174.780 295.600 175.420 ;
        RECT 4.000 173.420 295.600 174.780 ;
        RECT 4.000 172.700 296.000 173.420 ;
        RECT 4.400 172.020 296.000 172.700 ;
        RECT 4.400 170.700 295.600 172.020 ;
        RECT 4.000 170.020 295.600 170.700 ;
        RECT 4.000 168.620 296.000 170.020 ;
        RECT 4.400 166.620 295.600 168.620 ;
        RECT 4.000 165.220 296.000 166.620 ;
        RECT 4.000 164.540 295.600 165.220 ;
        RECT 4.400 163.220 295.600 164.540 ;
        RECT 4.400 162.540 296.000 163.220 ;
        RECT 4.000 161.140 296.000 162.540 ;
        RECT 4.000 160.460 295.600 161.140 ;
        RECT 4.400 159.140 295.600 160.460 ;
        RECT 4.400 158.460 296.000 159.140 ;
        RECT 4.000 157.740 296.000 158.460 ;
        RECT 4.000 156.380 295.600 157.740 ;
        RECT 4.400 155.740 295.600 156.380 ;
        RECT 4.400 154.380 296.000 155.740 ;
        RECT 4.000 154.340 296.000 154.380 ;
        RECT 4.000 152.340 295.600 154.340 ;
        RECT 4.000 152.300 296.000 152.340 ;
        RECT 4.400 150.940 296.000 152.300 ;
        RECT 4.400 150.300 295.600 150.940 ;
        RECT 4.000 148.940 295.600 150.300 ;
        RECT 4.000 148.220 296.000 148.940 ;
        RECT 4.400 147.540 296.000 148.220 ;
        RECT 4.400 146.220 295.600 147.540 ;
        RECT 4.000 145.540 295.600 146.220 ;
        RECT 4.000 144.140 296.000 145.540 ;
        RECT 4.400 142.140 295.600 144.140 ;
        RECT 4.000 140.740 296.000 142.140 ;
        RECT 4.400 138.740 295.600 140.740 ;
        RECT 4.000 137.340 296.000 138.740 ;
        RECT 4.000 136.660 295.600 137.340 ;
        RECT 4.400 135.340 295.600 136.660 ;
        RECT 4.400 134.660 296.000 135.340 ;
        RECT 4.000 133.940 296.000 134.660 ;
        RECT 4.000 132.580 295.600 133.940 ;
        RECT 4.400 131.940 295.600 132.580 ;
        RECT 4.400 130.580 296.000 131.940 ;
        RECT 4.000 130.540 296.000 130.580 ;
        RECT 4.000 128.540 295.600 130.540 ;
        RECT 4.000 128.500 296.000 128.540 ;
        RECT 4.400 127.140 296.000 128.500 ;
        RECT 4.400 126.500 295.600 127.140 ;
        RECT 4.000 125.140 295.600 126.500 ;
        RECT 4.000 124.420 296.000 125.140 ;
        RECT 4.400 123.740 296.000 124.420 ;
        RECT 4.400 122.420 295.600 123.740 ;
        RECT 4.000 121.740 295.600 122.420 ;
        RECT 4.000 120.340 296.000 121.740 ;
        RECT 4.400 119.660 296.000 120.340 ;
        RECT 4.400 118.340 295.600 119.660 ;
        RECT 4.000 117.660 295.600 118.340 ;
        RECT 4.000 116.260 296.000 117.660 ;
        RECT 4.400 114.260 295.600 116.260 ;
        RECT 4.000 112.860 296.000 114.260 ;
        RECT 4.000 112.180 295.600 112.860 ;
        RECT 4.400 110.860 295.600 112.180 ;
        RECT 4.400 110.180 296.000 110.860 ;
        RECT 4.000 109.460 296.000 110.180 ;
        RECT 4.000 108.100 295.600 109.460 ;
        RECT 4.400 107.460 295.600 108.100 ;
        RECT 4.400 106.100 296.000 107.460 ;
        RECT 4.000 106.060 296.000 106.100 ;
        RECT 4.000 104.060 295.600 106.060 ;
        RECT 4.000 104.020 296.000 104.060 ;
        RECT 4.400 102.660 296.000 104.020 ;
        RECT 4.400 102.020 295.600 102.660 ;
        RECT 4.000 100.660 295.600 102.020 ;
        RECT 4.000 99.940 296.000 100.660 ;
        RECT 4.400 99.260 296.000 99.940 ;
        RECT 4.400 97.940 295.600 99.260 ;
        RECT 4.000 97.260 295.600 97.940 ;
        RECT 4.000 95.860 296.000 97.260 ;
        RECT 4.400 93.860 295.600 95.860 ;
        RECT 4.000 92.460 296.000 93.860 ;
        RECT 4.000 91.780 295.600 92.460 ;
        RECT 4.400 90.460 295.600 91.780 ;
        RECT 4.400 89.780 296.000 90.460 ;
        RECT 4.000 89.060 296.000 89.780 ;
        RECT 4.000 87.700 295.600 89.060 ;
        RECT 4.400 87.060 295.600 87.700 ;
        RECT 4.400 85.700 296.000 87.060 ;
        RECT 4.000 85.660 296.000 85.700 ;
        RECT 4.000 83.660 295.600 85.660 ;
        RECT 4.000 83.620 296.000 83.660 ;
        RECT 4.400 81.620 296.000 83.620 ;
        RECT 4.000 81.580 296.000 81.620 ;
        RECT 4.000 79.580 295.600 81.580 ;
        RECT 4.000 79.540 296.000 79.580 ;
        RECT 4.400 78.180 296.000 79.540 ;
        RECT 4.400 77.540 295.600 78.180 ;
        RECT 4.000 76.180 295.600 77.540 ;
        RECT 4.000 75.460 296.000 76.180 ;
        RECT 4.400 74.780 296.000 75.460 ;
        RECT 4.400 73.460 295.600 74.780 ;
        RECT 4.000 72.780 295.600 73.460 ;
        RECT 4.000 71.380 296.000 72.780 ;
        RECT 4.400 69.380 295.600 71.380 ;
        RECT 4.000 67.980 296.000 69.380 ;
        RECT 4.000 67.300 295.600 67.980 ;
        RECT 4.400 65.980 295.600 67.300 ;
        RECT 4.400 65.300 296.000 65.980 ;
        RECT 4.000 64.580 296.000 65.300 ;
        RECT 4.000 63.220 295.600 64.580 ;
        RECT 4.400 62.580 295.600 63.220 ;
        RECT 4.400 61.220 296.000 62.580 ;
        RECT 4.000 61.180 296.000 61.220 ;
        RECT 4.000 59.180 295.600 61.180 ;
        RECT 4.000 59.140 296.000 59.180 ;
        RECT 4.400 57.780 296.000 59.140 ;
        RECT 4.400 57.140 295.600 57.780 ;
        RECT 4.000 55.780 295.600 57.140 ;
        RECT 4.000 55.060 296.000 55.780 ;
        RECT 4.400 54.380 296.000 55.060 ;
        RECT 4.400 53.060 295.600 54.380 ;
        RECT 4.000 52.380 295.600 53.060 ;
        RECT 4.000 50.980 296.000 52.380 ;
        RECT 4.400 48.980 295.600 50.980 ;
        RECT 4.000 47.580 296.000 48.980 ;
        RECT 4.000 46.900 295.600 47.580 ;
        RECT 4.400 45.580 295.600 46.900 ;
        RECT 4.400 44.900 296.000 45.580 ;
        RECT 4.000 44.180 296.000 44.900 ;
        RECT 4.000 42.820 295.600 44.180 ;
        RECT 4.400 42.180 295.600 42.820 ;
        RECT 4.400 40.820 296.000 42.180 ;
        RECT 4.000 40.100 296.000 40.820 ;
        RECT 4.000 38.740 295.600 40.100 ;
        RECT 4.400 38.100 295.600 38.740 ;
        RECT 4.400 36.740 296.000 38.100 ;
        RECT 4.000 36.700 296.000 36.740 ;
        RECT 4.000 34.700 295.600 36.700 ;
        RECT 4.000 34.660 296.000 34.700 ;
        RECT 4.400 33.300 296.000 34.660 ;
        RECT 4.400 32.660 295.600 33.300 ;
        RECT 4.000 31.300 295.600 32.660 ;
        RECT 4.000 30.580 296.000 31.300 ;
        RECT 4.400 29.900 296.000 30.580 ;
        RECT 4.400 28.580 295.600 29.900 ;
        RECT 4.000 27.900 295.600 28.580 ;
        RECT 4.000 26.500 296.000 27.900 ;
        RECT 4.400 24.500 295.600 26.500 ;
        RECT 4.000 23.100 296.000 24.500 ;
        RECT 4.000 22.420 295.600 23.100 ;
        RECT 4.400 21.100 295.600 22.420 ;
        RECT 4.400 20.420 296.000 21.100 ;
        RECT 4.000 19.700 296.000 20.420 ;
        RECT 4.000 18.340 295.600 19.700 ;
        RECT 4.400 17.700 295.600 18.340 ;
        RECT 4.400 16.340 296.000 17.700 ;
        RECT 4.000 16.300 296.000 16.340 ;
        RECT 4.000 14.300 295.600 16.300 ;
        RECT 4.000 14.260 296.000 14.300 ;
        RECT 4.400 12.900 296.000 14.260 ;
        RECT 4.400 12.260 295.600 12.900 ;
        RECT 4.000 10.900 295.600 12.260 ;
        RECT 4.000 10.180 296.000 10.900 ;
        RECT 4.400 9.500 296.000 10.180 ;
        RECT 4.400 8.180 295.600 9.500 ;
        RECT 4.000 7.500 295.600 8.180 ;
        RECT 4.000 6.100 296.000 7.500 ;
        RECT 4.400 4.100 295.600 6.100 ;
        RECT 4.000 2.700 296.000 4.100 ;
        RECT 4.400 2.555 295.600 2.700 ;
      LAYER met4 ;
        RECT 34.335 2.895 97.440 232.385 ;
        RECT 99.840 2.895 174.240 232.385 ;
        RECT 176.640 2.895 195.665 232.385 ;
  END
END wrapped_vgademo_on_fpga
END LIBRARY

