magic
tech sky130A
magscale 1 2
timestamp 1647824558
<< obsli1 >>
rect 1104 527 58880 57681
<< obsm1 >>
rect 658 496 59326 57996
<< metal2 >>
rect 634 59200 746 60000
rect 1922 59200 2034 60000
rect 3210 59200 3322 60000
rect 4498 59200 4610 60000
rect 5786 59200 5898 60000
rect 7074 59200 7186 60000
rect 8454 59200 8566 60000
rect 9742 59200 9854 60000
rect 11030 59200 11142 60000
rect 12318 59200 12430 60000
rect 13606 59200 13718 60000
rect 14894 59200 15006 60000
rect 16274 59200 16386 60000
rect 17562 59200 17674 60000
rect 18850 59200 18962 60000
rect 20138 59200 20250 60000
rect 21426 59200 21538 60000
rect 22714 59200 22826 60000
rect 24094 59200 24206 60000
rect 25382 59200 25494 60000
rect 26670 59200 26782 60000
rect 27958 59200 28070 60000
rect 29246 59200 29358 60000
rect 30626 59200 30738 60000
rect 31914 59200 32026 60000
rect 33202 59200 33314 60000
rect 34490 59200 34602 60000
rect 35778 59200 35890 60000
rect 37066 59200 37178 60000
rect 38446 59200 38558 60000
rect 39734 59200 39846 60000
rect 41022 59200 41134 60000
rect 42310 59200 42422 60000
rect 43598 59200 43710 60000
rect 44886 59200 44998 60000
rect 46266 59200 46378 60000
rect 47554 59200 47666 60000
rect 48842 59200 48954 60000
rect 50130 59200 50242 60000
rect 51418 59200 51530 60000
rect 52706 59200 52818 60000
rect 54086 59200 54198 60000
rect 55374 59200 55486 60000
rect 56662 59200 56774 60000
rect 57950 59200 58062 60000
rect 59238 59200 59350 60000
rect 2658 0 2770 800
rect 8086 0 8198 800
rect 13514 0 13626 800
rect 18942 0 19054 800
rect 24462 0 24574 800
rect 29890 0 30002 800
rect 35318 0 35430 800
rect 40746 0 40858 800
rect 46266 0 46378 800
rect 51694 0 51806 800
rect 57122 0 57234 800
<< obsm2 >>
rect 802 59144 1866 59537
rect 2090 59144 3154 59537
rect 3378 59144 4442 59537
rect 4666 59144 5730 59537
rect 5954 59144 7018 59537
rect 7242 59144 8398 59537
rect 8622 59144 9686 59537
rect 9910 59144 10974 59537
rect 11198 59144 12262 59537
rect 12486 59144 13550 59537
rect 13774 59144 14838 59537
rect 15062 59144 16218 59537
rect 16442 59144 17506 59537
rect 17730 59144 18794 59537
rect 19018 59144 20082 59537
rect 20306 59144 21370 59537
rect 21594 59144 22658 59537
rect 22882 59144 24038 59537
rect 24262 59144 25326 59537
rect 25550 59144 26614 59537
rect 26838 59144 27902 59537
rect 28126 59144 29190 59537
rect 29414 59144 30570 59537
rect 30794 59144 31858 59537
rect 32082 59144 33146 59537
rect 33370 59144 34434 59537
rect 34658 59144 35722 59537
rect 35946 59144 37010 59537
rect 37234 59144 38390 59537
rect 38614 59144 39678 59537
rect 39902 59144 40966 59537
rect 41190 59144 42254 59537
rect 42478 59144 43542 59537
rect 43766 59144 44830 59537
rect 45054 59144 46210 59537
rect 46434 59144 47498 59537
rect 47722 59144 48786 59537
rect 49010 59144 50074 59537
rect 50298 59144 51362 59537
rect 51586 59144 52650 59537
rect 52874 59144 54030 59537
rect 54254 59144 55318 59537
rect 55542 59144 56606 59537
rect 56830 59144 57894 59537
rect 58118 59144 59182 59537
rect 664 856 59320 59144
rect 664 496 2602 856
rect 2826 496 8030 856
rect 8254 496 13458 856
rect 13682 496 18886 856
rect 19110 496 24406 856
rect 24630 496 29834 856
rect 30058 496 35262 856
rect 35486 496 40690 856
rect 40914 496 46210 856
rect 46434 496 51638 856
rect 51862 496 57066 856
rect 57290 496 59320 856
<< metal3 >>
rect 0 59380 800 59620
rect 59200 59380 60000 59620
rect 0 58564 800 58804
rect 59200 58564 60000 58804
rect 0 57748 800 57988
rect 59200 57884 60000 58124
rect 0 56932 800 57172
rect 59200 57068 60000 57308
rect 0 56116 800 56356
rect 59200 56388 60000 56628
rect 0 55300 800 55540
rect 59200 55572 60000 55812
rect 59200 54892 60000 55132
rect 0 54484 800 54724
rect 59200 54076 60000 54316
rect 0 53668 800 53908
rect 59200 53396 60000 53636
rect 0 52988 800 53228
rect 59200 52580 60000 52820
rect 0 52172 800 52412
rect 59200 51900 60000 52140
rect 0 51356 800 51596
rect 59200 51084 60000 51324
rect 0 50540 800 50780
rect 59200 50404 60000 50644
rect 0 49724 800 49964
rect 59200 49588 60000 49828
rect 0 48908 800 49148
rect 59200 48908 60000 49148
rect 0 48092 800 48332
rect 59200 48092 60000 48332
rect 0 47276 800 47516
rect 59200 47412 60000 47652
rect 0 46596 800 46836
rect 59200 46596 60000 46836
rect 0 45780 800 46020
rect 59200 45916 60000 46156
rect 0 44964 800 45204
rect 59200 45100 60000 45340
rect 0 44148 800 44388
rect 59200 44420 60000 44660
rect 0 43332 800 43572
rect 59200 43604 60000 43844
rect 59200 42924 60000 43164
rect 0 42516 800 42756
rect 59200 42108 60000 42348
rect 0 41700 800 41940
rect 59200 41428 60000 41668
rect 0 40884 800 41124
rect 59200 40612 60000 40852
rect 0 40204 800 40444
rect 59200 39932 60000 40172
rect 0 39388 800 39628
rect 59200 39116 60000 39356
rect 0 38572 800 38812
rect 59200 38436 60000 38676
rect 0 37756 800 37996
rect 59200 37620 60000 37860
rect 0 36940 800 37180
rect 59200 36940 60000 37180
rect 0 36124 800 36364
rect 59200 36124 60000 36364
rect 0 35308 800 35548
rect 59200 35444 60000 35684
rect 0 34492 800 34732
rect 59200 34628 60000 34868
rect 0 33676 800 33916
rect 59200 33948 60000 34188
rect 0 32996 800 33236
rect 59200 33132 60000 33372
rect 0 32180 800 32420
rect 59200 32452 60000 32692
rect 0 31364 800 31604
rect 59200 31636 60000 31876
rect 59200 30956 60000 31196
rect 0 30548 800 30788
rect 59200 30140 60000 30380
rect 0 29732 800 29972
rect 59200 29324 60000 29564
rect 0 28916 800 29156
rect 59200 28644 60000 28884
rect 0 28100 800 28340
rect 59200 27828 60000 28068
rect 0 27284 800 27524
rect 59200 27148 60000 27388
rect 0 26604 800 26844
rect 59200 26332 60000 26572
rect 0 25788 800 26028
rect 59200 25652 60000 25892
rect 0 24972 800 25212
rect 59200 24836 60000 25076
rect 0 24156 800 24396
rect 59200 24156 60000 24396
rect 0 23340 800 23580
rect 59200 23340 60000 23580
rect 0 22524 800 22764
rect 59200 22660 60000 22900
rect 0 21708 800 21948
rect 59200 21844 60000 22084
rect 0 20892 800 21132
rect 59200 21164 60000 21404
rect 0 20212 800 20452
rect 59200 20348 60000 20588
rect 0 19396 800 19636
rect 59200 19668 60000 19908
rect 0 18580 800 18820
rect 59200 18852 60000 19092
rect 59200 18172 60000 18412
rect 0 17764 800 18004
rect 59200 17356 60000 17596
rect 0 16948 800 17188
rect 59200 16676 60000 16916
rect 0 16132 800 16372
rect 59200 15860 60000 16100
rect 0 15316 800 15556
rect 59200 15180 60000 15420
rect 0 14500 800 14740
rect 59200 14364 60000 14604
rect 0 13684 800 13924
rect 59200 13684 60000 13924
rect 0 13004 800 13244
rect 59200 12868 60000 13108
rect 0 12188 800 12428
rect 59200 12188 60000 12428
rect 0 11372 800 11612
rect 59200 11372 60000 11612
rect 0 10556 800 10796
rect 59200 10692 60000 10932
rect 0 9740 800 9980
rect 59200 9876 60000 10116
rect 0 8924 800 9164
rect 59200 9196 60000 9436
rect 0 8108 800 8348
rect 59200 8380 60000 8620
rect 59200 7700 60000 7940
rect 0 7292 800 7532
rect 0 6612 800 6852
rect 59200 6884 60000 7124
rect 59200 6204 60000 6444
rect 0 5796 800 6036
rect 59200 5388 60000 5628
rect 0 4980 800 5220
rect 59200 4708 60000 4948
rect 0 4164 800 4404
rect 59200 3892 60000 4132
rect 0 3348 800 3588
rect 59200 3212 60000 3452
rect 0 2532 800 2772
rect 59200 2396 60000 2636
rect 0 1716 800 1956
rect 59200 1716 60000 1956
rect 0 900 800 1140
rect 59200 900 60000 1140
rect 0 220 800 460
rect 59200 220 60000 460
<< obsm3 >>
rect 880 59300 59120 59533
rect 800 58884 59200 59300
rect 880 58484 59120 58884
rect 800 58204 59200 58484
rect 800 58068 59120 58204
rect 880 57804 59120 58068
rect 880 57668 59200 57804
rect 800 57388 59200 57668
rect 800 57252 59120 57388
rect 880 56988 59120 57252
rect 880 56852 59200 56988
rect 800 56708 59200 56852
rect 800 56436 59120 56708
rect 880 56308 59120 56436
rect 880 56036 59200 56308
rect 800 55892 59200 56036
rect 800 55620 59120 55892
rect 880 55492 59120 55620
rect 880 55220 59200 55492
rect 800 55212 59200 55220
rect 800 54812 59120 55212
rect 800 54804 59200 54812
rect 880 54404 59200 54804
rect 800 54396 59200 54404
rect 800 53996 59120 54396
rect 800 53988 59200 53996
rect 880 53716 59200 53988
rect 880 53588 59120 53716
rect 800 53316 59120 53588
rect 800 53308 59200 53316
rect 880 52908 59200 53308
rect 800 52900 59200 52908
rect 800 52500 59120 52900
rect 800 52492 59200 52500
rect 880 52220 59200 52492
rect 880 52092 59120 52220
rect 800 51820 59120 52092
rect 800 51676 59200 51820
rect 880 51404 59200 51676
rect 880 51276 59120 51404
rect 800 51004 59120 51276
rect 800 50860 59200 51004
rect 880 50724 59200 50860
rect 880 50460 59120 50724
rect 800 50324 59120 50460
rect 800 50044 59200 50324
rect 880 49908 59200 50044
rect 880 49644 59120 49908
rect 800 49508 59120 49644
rect 800 49228 59200 49508
rect 880 48828 59120 49228
rect 800 48412 59200 48828
rect 880 48012 59120 48412
rect 800 47732 59200 48012
rect 800 47596 59120 47732
rect 880 47332 59120 47596
rect 880 47196 59200 47332
rect 800 46916 59200 47196
rect 880 46516 59120 46916
rect 800 46236 59200 46516
rect 800 46100 59120 46236
rect 880 45836 59120 46100
rect 880 45700 59200 45836
rect 800 45420 59200 45700
rect 800 45284 59120 45420
rect 880 45020 59120 45284
rect 880 44884 59200 45020
rect 800 44740 59200 44884
rect 800 44468 59120 44740
rect 880 44340 59120 44468
rect 880 44068 59200 44340
rect 800 43924 59200 44068
rect 800 43652 59120 43924
rect 880 43524 59120 43652
rect 880 43252 59200 43524
rect 800 43244 59200 43252
rect 800 42844 59120 43244
rect 800 42836 59200 42844
rect 880 42436 59200 42836
rect 800 42428 59200 42436
rect 800 42028 59120 42428
rect 800 42020 59200 42028
rect 880 41748 59200 42020
rect 880 41620 59120 41748
rect 800 41348 59120 41620
rect 800 41204 59200 41348
rect 880 40932 59200 41204
rect 880 40804 59120 40932
rect 800 40532 59120 40804
rect 800 40524 59200 40532
rect 880 40252 59200 40524
rect 880 40124 59120 40252
rect 800 39852 59120 40124
rect 800 39708 59200 39852
rect 880 39436 59200 39708
rect 880 39308 59120 39436
rect 800 39036 59120 39308
rect 800 38892 59200 39036
rect 880 38756 59200 38892
rect 880 38492 59120 38756
rect 800 38356 59120 38492
rect 800 38076 59200 38356
rect 880 37940 59200 38076
rect 880 37676 59120 37940
rect 800 37540 59120 37676
rect 800 37260 59200 37540
rect 880 36860 59120 37260
rect 800 36444 59200 36860
rect 880 36044 59120 36444
rect 800 35764 59200 36044
rect 800 35628 59120 35764
rect 880 35364 59120 35628
rect 880 35228 59200 35364
rect 800 34948 59200 35228
rect 800 34812 59120 34948
rect 880 34548 59120 34812
rect 880 34412 59200 34548
rect 800 34268 59200 34412
rect 800 33996 59120 34268
rect 880 33868 59120 33996
rect 880 33596 59200 33868
rect 800 33452 59200 33596
rect 800 33316 59120 33452
rect 880 33052 59120 33316
rect 880 32916 59200 33052
rect 800 32772 59200 32916
rect 800 32500 59120 32772
rect 880 32372 59120 32500
rect 880 32100 59200 32372
rect 800 31956 59200 32100
rect 800 31684 59120 31956
rect 880 31556 59120 31684
rect 880 31284 59200 31556
rect 800 31276 59200 31284
rect 800 30876 59120 31276
rect 800 30868 59200 30876
rect 880 30468 59200 30868
rect 800 30460 59200 30468
rect 800 30060 59120 30460
rect 800 30052 59200 30060
rect 880 29652 59200 30052
rect 800 29644 59200 29652
rect 800 29244 59120 29644
rect 800 29236 59200 29244
rect 880 28964 59200 29236
rect 880 28836 59120 28964
rect 800 28564 59120 28836
rect 800 28420 59200 28564
rect 880 28148 59200 28420
rect 880 28020 59120 28148
rect 800 27748 59120 28020
rect 800 27604 59200 27748
rect 880 27468 59200 27604
rect 880 27204 59120 27468
rect 800 27068 59120 27204
rect 800 26924 59200 27068
rect 880 26652 59200 26924
rect 880 26524 59120 26652
rect 800 26252 59120 26524
rect 800 26108 59200 26252
rect 880 25972 59200 26108
rect 880 25708 59120 25972
rect 800 25572 59120 25708
rect 800 25292 59200 25572
rect 880 25156 59200 25292
rect 880 24892 59120 25156
rect 800 24756 59120 24892
rect 800 24476 59200 24756
rect 880 24076 59120 24476
rect 800 23660 59200 24076
rect 880 23260 59120 23660
rect 800 22980 59200 23260
rect 800 22844 59120 22980
rect 880 22580 59120 22844
rect 880 22444 59200 22580
rect 800 22164 59200 22444
rect 800 22028 59120 22164
rect 880 21764 59120 22028
rect 880 21628 59200 21764
rect 800 21484 59200 21628
rect 800 21212 59120 21484
rect 880 21084 59120 21212
rect 880 20812 59200 21084
rect 800 20668 59200 20812
rect 800 20532 59120 20668
rect 880 20268 59120 20532
rect 880 20132 59200 20268
rect 800 19988 59200 20132
rect 800 19716 59120 19988
rect 880 19588 59120 19716
rect 880 19316 59200 19588
rect 800 19172 59200 19316
rect 800 18900 59120 19172
rect 880 18772 59120 18900
rect 880 18500 59200 18772
rect 800 18492 59200 18500
rect 800 18092 59120 18492
rect 800 18084 59200 18092
rect 880 17684 59200 18084
rect 800 17676 59200 17684
rect 800 17276 59120 17676
rect 800 17268 59200 17276
rect 880 16996 59200 17268
rect 880 16868 59120 16996
rect 800 16596 59120 16868
rect 800 16452 59200 16596
rect 880 16180 59200 16452
rect 880 16052 59120 16180
rect 800 15780 59120 16052
rect 800 15636 59200 15780
rect 880 15500 59200 15636
rect 880 15236 59120 15500
rect 800 15100 59120 15236
rect 800 14820 59200 15100
rect 880 14684 59200 14820
rect 880 14420 59120 14684
rect 800 14284 59120 14420
rect 800 14004 59200 14284
rect 880 13604 59120 14004
rect 800 13324 59200 13604
rect 880 13188 59200 13324
rect 880 12924 59120 13188
rect 800 12788 59120 12924
rect 800 12508 59200 12788
rect 880 12108 59120 12508
rect 800 11692 59200 12108
rect 880 11292 59120 11692
rect 800 11012 59200 11292
rect 800 10876 59120 11012
rect 880 10612 59120 10876
rect 880 10476 59200 10612
rect 800 10196 59200 10476
rect 800 10060 59120 10196
rect 880 9796 59120 10060
rect 880 9660 59200 9796
rect 800 9516 59200 9660
rect 800 9244 59120 9516
rect 880 9116 59120 9244
rect 880 8844 59200 9116
rect 800 8700 59200 8844
rect 800 8428 59120 8700
rect 880 8300 59120 8428
rect 880 8028 59200 8300
rect 800 8020 59200 8028
rect 800 7620 59120 8020
rect 800 7612 59200 7620
rect 880 7212 59200 7612
rect 800 7204 59200 7212
rect 800 6932 59120 7204
rect 880 6804 59120 6932
rect 880 6532 59200 6804
rect 800 6524 59200 6532
rect 800 6124 59120 6524
rect 800 6116 59200 6124
rect 880 5716 59200 6116
rect 800 5708 59200 5716
rect 800 5308 59120 5708
rect 800 5300 59200 5308
rect 880 5028 59200 5300
rect 880 4900 59120 5028
rect 800 4628 59120 4900
rect 800 4484 59200 4628
rect 880 4212 59200 4484
rect 880 4084 59120 4212
rect 800 3812 59120 4084
rect 800 3668 59200 3812
rect 880 3532 59200 3668
rect 880 3268 59120 3532
rect 800 3132 59120 3268
rect 800 2852 59200 3132
rect 880 2716 59200 2852
rect 880 2452 59120 2716
rect 800 2316 59120 2452
rect 800 2036 59200 2316
rect 880 1636 59120 2036
rect 800 1220 59200 1636
rect 880 820 59120 1220
rect 800 540 59200 820
rect 880 511 59120 540
<< metal4 >>
rect 4208 496 4528 57712
rect 19568 496 19888 57712
rect 34928 496 35248 57712
rect 50288 496 50608 57712
<< obsm4 >>
rect 4659 1395 19488 54501
rect 19968 1395 34848 54501
rect 35328 1395 49989 54501
<< labels >>
rlabel metal2 s 634 59200 746 60000 6 active
port 1 nsew signal input
rlabel metal2 s 3210 59200 3322 60000 6 io_in[0]
port 2 nsew signal input
rlabel metal2 s 16274 59200 16386 60000 6 io_in[10]
port 3 nsew signal input
rlabel metal2 s 17562 59200 17674 60000 6 io_in[11]
port 4 nsew signal input
rlabel metal2 s 18850 59200 18962 60000 6 io_in[12]
port 5 nsew signal input
rlabel metal2 s 20138 59200 20250 60000 6 io_in[13]
port 6 nsew signal input
rlabel metal2 s 21426 59200 21538 60000 6 io_in[14]
port 7 nsew signal input
rlabel metal2 s 22714 59200 22826 60000 6 io_in[15]
port 8 nsew signal input
rlabel metal2 s 24094 59200 24206 60000 6 io_in[16]
port 9 nsew signal input
rlabel metal2 s 25382 59200 25494 60000 6 io_in[17]
port 10 nsew signal input
rlabel metal2 s 26670 59200 26782 60000 6 io_in[18]
port 11 nsew signal input
rlabel metal2 s 27958 59200 28070 60000 6 io_in[19]
port 12 nsew signal input
rlabel metal2 s 4498 59200 4610 60000 6 io_in[1]
port 13 nsew signal input
rlabel metal2 s 29246 59200 29358 60000 6 io_in[20]
port 14 nsew signal input
rlabel metal2 s 30626 59200 30738 60000 6 io_in[21]
port 15 nsew signal input
rlabel metal2 s 31914 59200 32026 60000 6 io_in[22]
port 16 nsew signal input
rlabel metal2 s 33202 59200 33314 60000 6 io_in[23]
port 17 nsew signal input
rlabel metal2 s 34490 59200 34602 60000 6 io_in[24]
port 18 nsew signal input
rlabel metal2 s 35778 59200 35890 60000 6 io_in[25]
port 19 nsew signal input
rlabel metal2 s 37066 59200 37178 60000 6 io_in[26]
port 20 nsew signal input
rlabel metal2 s 38446 59200 38558 60000 6 io_in[27]
port 21 nsew signal input
rlabel metal2 s 39734 59200 39846 60000 6 io_in[28]
port 22 nsew signal input
rlabel metal2 s 41022 59200 41134 60000 6 io_in[29]
port 23 nsew signal input
rlabel metal2 s 5786 59200 5898 60000 6 io_in[2]
port 24 nsew signal input
rlabel metal2 s 42310 59200 42422 60000 6 io_in[30]
port 25 nsew signal input
rlabel metal2 s 43598 59200 43710 60000 6 io_in[31]
port 26 nsew signal input
rlabel metal2 s 44886 59200 44998 60000 6 io_in[32]
port 27 nsew signal input
rlabel metal2 s 46266 59200 46378 60000 6 io_in[33]
port 28 nsew signal input
rlabel metal2 s 47554 59200 47666 60000 6 io_in[34]
port 29 nsew signal input
rlabel metal2 s 48842 59200 48954 60000 6 io_in[35]
port 30 nsew signal input
rlabel metal2 s 50130 59200 50242 60000 6 io_in[36]
port 31 nsew signal input
rlabel metal2 s 51418 59200 51530 60000 6 io_in[37]
port 32 nsew signal input
rlabel metal2 s 7074 59200 7186 60000 6 io_in[3]
port 33 nsew signal input
rlabel metal2 s 8454 59200 8566 60000 6 io_in[4]
port 34 nsew signal input
rlabel metal2 s 9742 59200 9854 60000 6 io_in[5]
port 35 nsew signal input
rlabel metal2 s 11030 59200 11142 60000 6 io_in[6]
port 36 nsew signal input
rlabel metal2 s 12318 59200 12430 60000 6 io_in[7]
port 37 nsew signal input
rlabel metal2 s 13606 59200 13718 60000 6 io_in[8]
port 38 nsew signal input
rlabel metal2 s 14894 59200 15006 60000 6 io_in[9]
port 39 nsew signal input
rlabel metal3 s 59200 24156 60000 24396 6 io_oeb[0]
port 40 nsew signal output
rlabel metal3 s 59200 31636 60000 31876 6 io_oeb[10]
port 41 nsew signal output
rlabel metal3 s 59200 32452 60000 32692 6 io_oeb[11]
port 42 nsew signal output
rlabel metal3 s 59200 33132 60000 33372 6 io_oeb[12]
port 43 nsew signal output
rlabel metal3 s 59200 33948 60000 34188 6 io_oeb[13]
port 44 nsew signal output
rlabel metal3 s 59200 34628 60000 34868 6 io_oeb[14]
port 45 nsew signal output
rlabel metal3 s 59200 35444 60000 35684 6 io_oeb[15]
port 46 nsew signal output
rlabel metal3 s 59200 36124 60000 36364 6 io_oeb[16]
port 47 nsew signal output
rlabel metal3 s 59200 36940 60000 37180 6 io_oeb[17]
port 48 nsew signal output
rlabel metal3 s 59200 37620 60000 37860 6 io_oeb[18]
port 49 nsew signal output
rlabel metal3 s 59200 38436 60000 38676 6 io_oeb[19]
port 50 nsew signal output
rlabel metal3 s 59200 24836 60000 25076 6 io_oeb[1]
port 51 nsew signal output
rlabel metal3 s 59200 39116 60000 39356 6 io_oeb[20]
port 52 nsew signal output
rlabel metal3 s 59200 39932 60000 40172 6 io_oeb[21]
port 53 nsew signal output
rlabel metal3 s 59200 40612 60000 40852 6 io_oeb[22]
port 54 nsew signal output
rlabel metal3 s 59200 41428 60000 41668 6 io_oeb[23]
port 55 nsew signal output
rlabel metal3 s 59200 42108 60000 42348 6 io_oeb[24]
port 56 nsew signal output
rlabel metal3 s 59200 42924 60000 43164 6 io_oeb[25]
port 57 nsew signal output
rlabel metal3 s 59200 43604 60000 43844 6 io_oeb[26]
port 58 nsew signal output
rlabel metal3 s 59200 44420 60000 44660 6 io_oeb[27]
port 59 nsew signal output
rlabel metal3 s 59200 45100 60000 45340 6 io_oeb[28]
port 60 nsew signal output
rlabel metal3 s 59200 45916 60000 46156 6 io_oeb[29]
port 61 nsew signal output
rlabel metal3 s 59200 25652 60000 25892 6 io_oeb[2]
port 62 nsew signal output
rlabel metal3 s 59200 46596 60000 46836 6 io_oeb[30]
port 63 nsew signal output
rlabel metal3 s 59200 47412 60000 47652 6 io_oeb[31]
port 64 nsew signal output
rlabel metal3 s 59200 48092 60000 48332 6 io_oeb[32]
port 65 nsew signal output
rlabel metal3 s 59200 48908 60000 49148 6 io_oeb[33]
port 66 nsew signal output
rlabel metal3 s 59200 49588 60000 49828 6 io_oeb[34]
port 67 nsew signal output
rlabel metal3 s 59200 50404 60000 50644 6 io_oeb[35]
port 68 nsew signal output
rlabel metal3 s 59200 51084 60000 51324 6 io_oeb[36]
port 69 nsew signal output
rlabel metal3 s 59200 51900 60000 52140 6 io_oeb[37]
port 70 nsew signal output
rlabel metal3 s 59200 26332 60000 26572 6 io_oeb[3]
port 71 nsew signal output
rlabel metal3 s 59200 27148 60000 27388 6 io_oeb[4]
port 72 nsew signal output
rlabel metal3 s 59200 27828 60000 28068 6 io_oeb[5]
port 73 nsew signal output
rlabel metal3 s 59200 28644 60000 28884 6 io_oeb[6]
port 74 nsew signal output
rlabel metal3 s 59200 29324 60000 29564 6 io_oeb[7]
port 75 nsew signal output
rlabel metal3 s 59200 30140 60000 30380 6 io_oeb[8]
port 76 nsew signal output
rlabel metal3 s 59200 30956 60000 31196 6 io_oeb[9]
port 77 nsew signal output
rlabel metal3 s 0 51356 800 51596 6 io_out[0]
port 78 nsew signal output
rlabel metal3 s 59200 54076 60000 54316 6 io_out[10]
port 79 nsew signal output
rlabel metal2 s 18942 0 19054 800 6 io_out[11]
port 80 nsew signal output
rlabel metal2 s 55374 59200 55486 60000 6 io_out[12]
port 81 nsew signal output
rlabel metal3 s 0 53668 800 53908 6 io_out[13]
port 82 nsew signal output
rlabel metal2 s 24462 0 24574 800 6 io_out[14]
port 83 nsew signal output
rlabel metal3 s 59200 54892 60000 55132 6 io_out[15]
port 84 nsew signal output
rlabel metal2 s 29890 0 30002 800 6 io_out[16]
port 85 nsew signal output
rlabel metal2 s 35318 0 35430 800 6 io_out[17]
port 86 nsew signal output
rlabel metal2 s 40746 0 40858 800 6 io_out[18]
port 87 nsew signal output
rlabel metal2 s 46266 0 46378 800 6 io_out[19]
port 88 nsew signal output
rlabel metal2 s 2658 0 2770 800 6 io_out[1]
port 89 nsew signal output
rlabel metal3 s 0 54484 800 54724 6 io_out[20]
port 90 nsew signal output
rlabel metal2 s 51694 0 51806 800 6 io_out[21]
port 91 nsew signal output
rlabel metal3 s 0 55300 800 55540 6 io_out[22]
port 92 nsew signal output
rlabel metal3 s 59200 55572 60000 55812 6 io_out[23]
port 93 nsew signal output
rlabel metal2 s 57122 0 57234 800 6 io_out[24]
port 94 nsew signal output
rlabel metal3 s 0 56116 800 56356 6 io_out[25]
port 95 nsew signal output
rlabel metal3 s 0 56932 800 57172 6 io_out[26]
port 96 nsew signal output
rlabel metal3 s 59200 56388 60000 56628 6 io_out[27]
port 97 nsew signal output
rlabel metal3 s 0 57748 800 57988 6 io_out[28]
port 98 nsew signal output
rlabel metal3 s 59200 57068 60000 57308 6 io_out[29]
port 99 nsew signal output
rlabel metal3 s 59200 52580 60000 52820 6 io_out[2]
port 100 nsew signal output
rlabel metal2 s 56662 59200 56774 60000 6 io_out[30]
port 101 nsew signal output
rlabel metal3 s 59200 57884 60000 58124 6 io_out[31]
port 102 nsew signal output
rlabel metal3 s 0 58564 800 58804 6 io_out[32]
port 103 nsew signal output
rlabel metal3 s 0 59380 800 59620 6 io_out[33]
port 104 nsew signal output
rlabel metal2 s 57950 59200 58062 60000 6 io_out[34]
port 105 nsew signal output
rlabel metal3 s 59200 58564 60000 58804 6 io_out[35]
port 106 nsew signal output
rlabel metal3 s 59200 59380 60000 59620 6 io_out[36]
port 107 nsew signal output
rlabel metal2 s 59238 59200 59350 60000 6 io_out[37]
port 108 nsew signal output
rlabel metal2 s 52706 59200 52818 60000 6 io_out[3]
port 109 nsew signal output
rlabel metal3 s 0 52172 800 52412 6 io_out[4]
port 110 nsew signal output
rlabel metal3 s 0 52988 800 53228 6 io_out[5]
port 111 nsew signal output
rlabel metal2 s 54086 59200 54198 60000 6 io_out[6]
port 112 nsew signal output
rlabel metal3 s 59200 53396 60000 53636 6 io_out[7]
port 113 nsew signal output
rlabel metal2 s 8086 0 8198 800 6 io_out[8]
port 114 nsew signal output
rlabel metal2 s 13514 0 13626 800 6 io_out[9]
port 115 nsew signal output
rlabel metal3 s 0 220 800 460 6 la1_data_in[0]
port 116 nsew signal input
rlabel metal3 s 0 8108 800 8348 6 la1_data_in[10]
port 117 nsew signal input
rlabel metal3 s 0 8924 800 9164 6 la1_data_in[11]
port 118 nsew signal input
rlabel metal3 s 0 9740 800 9980 6 la1_data_in[12]
port 119 nsew signal input
rlabel metal3 s 0 10556 800 10796 6 la1_data_in[13]
port 120 nsew signal input
rlabel metal3 s 0 11372 800 11612 6 la1_data_in[14]
port 121 nsew signal input
rlabel metal3 s 0 12188 800 12428 6 la1_data_in[15]
port 122 nsew signal input
rlabel metal3 s 0 13004 800 13244 6 la1_data_in[16]
port 123 nsew signal input
rlabel metal3 s 0 13684 800 13924 6 la1_data_in[17]
port 124 nsew signal input
rlabel metal3 s 0 14500 800 14740 6 la1_data_in[18]
port 125 nsew signal input
rlabel metal3 s 0 15316 800 15556 6 la1_data_in[19]
port 126 nsew signal input
rlabel metal3 s 0 900 800 1140 6 la1_data_in[1]
port 127 nsew signal input
rlabel metal3 s 0 16132 800 16372 6 la1_data_in[20]
port 128 nsew signal input
rlabel metal3 s 0 16948 800 17188 6 la1_data_in[21]
port 129 nsew signal input
rlabel metal3 s 0 17764 800 18004 6 la1_data_in[22]
port 130 nsew signal input
rlabel metal3 s 0 18580 800 18820 6 la1_data_in[23]
port 131 nsew signal input
rlabel metal3 s 0 19396 800 19636 6 la1_data_in[24]
port 132 nsew signal input
rlabel metal3 s 0 20212 800 20452 6 la1_data_in[25]
port 133 nsew signal input
rlabel metal3 s 0 20892 800 21132 6 la1_data_in[26]
port 134 nsew signal input
rlabel metal3 s 0 21708 800 21948 6 la1_data_in[27]
port 135 nsew signal input
rlabel metal3 s 0 22524 800 22764 6 la1_data_in[28]
port 136 nsew signal input
rlabel metal3 s 0 23340 800 23580 6 la1_data_in[29]
port 137 nsew signal input
rlabel metal3 s 0 1716 800 1956 6 la1_data_in[2]
port 138 nsew signal input
rlabel metal3 s 0 24156 800 24396 6 la1_data_in[30]
port 139 nsew signal input
rlabel metal3 s 0 24972 800 25212 6 la1_data_in[31]
port 140 nsew signal input
rlabel metal3 s 0 2532 800 2772 6 la1_data_in[3]
port 141 nsew signal input
rlabel metal3 s 0 3348 800 3588 6 la1_data_in[4]
port 142 nsew signal input
rlabel metal3 s 0 4164 800 4404 6 la1_data_in[5]
port 143 nsew signal input
rlabel metal3 s 0 4980 800 5220 6 la1_data_in[6]
port 144 nsew signal input
rlabel metal3 s 0 5796 800 6036 6 la1_data_in[7]
port 145 nsew signal input
rlabel metal3 s 0 6612 800 6852 6 la1_data_in[8]
port 146 nsew signal input
rlabel metal3 s 0 7292 800 7532 6 la1_data_in[9]
port 147 nsew signal input
rlabel metal3 s 0 25788 800 26028 6 la1_data_out[0]
port 148 nsew signal output
rlabel metal3 s 0 33676 800 33916 6 la1_data_out[10]
port 149 nsew signal output
rlabel metal3 s 0 34492 800 34732 6 la1_data_out[11]
port 150 nsew signal output
rlabel metal3 s 0 35308 800 35548 6 la1_data_out[12]
port 151 nsew signal output
rlabel metal3 s 0 36124 800 36364 6 la1_data_out[13]
port 152 nsew signal output
rlabel metal3 s 0 36940 800 37180 6 la1_data_out[14]
port 153 nsew signal output
rlabel metal3 s 0 37756 800 37996 6 la1_data_out[15]
port 154 nsew signal output
rlabel metal3 s 0 38572 800 38812 6 la1_data_out[16]
port 155 nsew signal output
rlabel metal3 s 0 39388 800 39628 6 la1_data_out[17]
port 156 nsew signal output
rlabel metal3 s 0 40204 800 40444 6 la1_data_out[18]
port 157 nsew signal output
rlabel metal3 s 0 40884 800 41124 6 la1_data_out[19]
port 158 nsew signal output
rlabel metal3 s 0 26604 800 26844 6 la1_data_out[1]
port 159 nsew signal output
rlabel metal3 s 0 41700 800 41940 6 la1_data_out[20]
port 160 nsew signal output
rlabel metal3 s 0 42516 800 42756 6 la1_data_out[21]
port 161 nsew signal output
rlabel metal3 s 0 43332 800 43572 6 la1_data_out[22]
port 162 nsew signal output
rlabel metal3 s 0 44148 800 44388 6 la1_data_out[23]
port 163 nsew signal output
rlabel metal3 s 0 44964 800 45204 6 la1_data_out[24]
port 164 nsew signal output
rlabel metal3 s 0 45780 800 46020 6 la1_data_out[25]
port 165 nsew signal output
rlabel metal3 s 0 46596 800 46836 6 la1_data_out[26]
port 166 nsew signal output
rlabel metal3 s 0 47276 800 47516 6 la1_data_out[27]
port 167 nsew signal output
rlabel metal3 s 0 48092 800 48332 6 la1_data_out[28]
port 168 nsew signal output
rlabel metal3 s 0 48908 800 49148 6 la1_data_out[29]
port 169 nsew signal output
rlabel metal3 s 0 27284 800 27524 6 la1_data_out[2]
port 170 nsew signal output
rlabel metal3 s 0 49724 800 49964 6 la1_data_out[30]
port 171 nsew signal output
rlabel metal3 s 0 50540 800 50780 6 la1_data_out[31]
port 172 nsew signal output
rlabel metal3 s 0 28100 800 28340 6 la1_data_out[3]
port 173 nsew signal output
rlabel metal3 s 0 28916 800 29156 6 la1_data_out[4]
port 174 nsew signal output
rlabel metal3 s 0 29732 800 29972 6 la1_data_out[5]
port 175 nsew signal output
rlabel metal3 s 0 30548 800 30788 6 la1_data_out[6]
port 176 nsew signal output
rlabel metal3 s 0 31364 800 31604 6 la1_data_out[7]
port 177 nsew signal output
rlabel metal3 s 0 32180 800 32420 6 la1_data_out[8]
port 178 nsew signal output
rlabel metal3 s 0 32996 800 33236 6 la1_data_out[9]
port 179 nsew signal output
rlabel metal3 s 59200 220 60000 460 6 la1_oenb[0]
port 180 nsew signal input
rlabel metal3 s 59200 7700 60000 7940 6 la1_oenb[10]
port 181 nsew signal input
rlabel metal3 s 59200 8380 60000 8620 6 la1_oenb[11]
port 182 nsew signal input
rlabel metal3 s 59200 9196 60000 9436 6 la1_oenb[12]
port 183 nsew signal input
rlabel metal3 s 59200 9876 60000 10116 6 la1_oenb[13]
port 184 nsew signal input
rlabel metal3 s 59200 10692 60000 10932 6 la1_oenb[14]
port 185 nsew signal input
rlabel metal3 s 59200 11372 60000 11612 6 la1_oenb[15]
port 186 nsew signal input
rlabel metal3 s 59200 12188 60000 12428 6 la1_oenb[16]
port 187 nsew signal input
rlabel metal3 s 59200 12868 60000 13108 6 la1_oenb[17]
port 188 nsew signal input
rlabel metal3 s 59200 13684 60000 13924 6 la1_oenb[18]
port 189 nsew signal input
rlabel metal3 s 59200 14364 60000 14604 6 la1_oenb[19]
port 190 nsew signal input
rlabel metal3 s 59200 900 60000 1140 6 la1_oenb[1]
port 191 nsew signal input
rlabel metal3 s 59200 15180 60000 15420 6 la1_oenb[20]
port 192 nsew signal input
rlabel metal3 s 59200 15860 60000 16100 6 la1_oenb[21]
port 193 nsew signal input
rlabel metal3 s 59200 16676 60000 16916 6 la1_oenb[22]
port 194 nsew signal input
rlabel metal3 s 59200 17356 60000 17596 6 la1_oenb[23]
port 195 nsew signal input
rlabel metal3 s 59200 18172 60000 18412 6 la1_oenb[24]
port 196 nsew signal input
rlabel metal3 s 59200 18852 60000 19092 6 la1_oenb[25]
port 197 nsew signal input
rlabel metal3 s 59200 19668 60000 19908 6 la1_oenb[26]
port 198 nsew signal input
rlabel metal3 s 59200 20348 60000 20588 6 la1_oenb[27]
port 199 nsew signal input
rlabel metal3 s 59200 21164 60000 21404 6 la1_oenb[28]
port 200 nsew signal input
rlabel metal3 s 59200 21844 60000 22084 6 la1_oenb[29]
port 201 nsew signal input
rlabel metal3 s 59200 1716 60000 1956 6 la1_oenb[2]
port 202 nsew signal input
rlabel metal3 s 59200 22660 60000 22900 6 la1_oenb[30]
port 203 nsew signal input
rlabel metal3 s 59200 23340 60000 23580 6 la1_oenb[31]
port 204 nsew signal input
rlabel metal3 s 59200 2396 60000 2636 6 la1_oenb[3]
port 205 nsew signal input
rlabel metal3 s 59200 3212 60000 3452 6 la1_oenb[4]
port 206 nsew signal input
rlabel metal3 s 59200 3892 60000 4132 6 la1_oenb[5]
port 207 nsew signal input
rlabel metal3 s 59200 4708 60000 4948 6 la1_oenb[6]
port 208 nsew signal input
rlabel metal3 s 59200 5388 60000 5628 6 la1_oenb[7]
port 209 nsew signal input
rlabel metal3 s 59200 6204 60000 6444 6 la1_oenb[8]
port 210 nsew signal input
rlabel metal3 s 59200 6884 60000 7124 6 la1_oenb[9]
port 211 nsew signal input
rlabel metal4 s 4208 496 4528 57712 6 vccd1
port 212 nsew power input
rlabel metal4 s 34928 496 35248 57712 6 vccd1
port 212 nsew power input
rlabel metal4 s 19568 496 19888 57712 6 vssd1
port 213 nsew ground input
rlabel metal4 s 50288 496 50608 57712 6 vssd1
port 213 nsew ground input
rlabel metal2 s 1922 59200 2034 60000 6 wb_clk_i
port 214 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 60000 60000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 12736066
string GDS_FILE /openlane/designs/wrapped-vgademo-on-fpga/runs/RUN_2022.03.21_00.58.11/results/finishing/wrapped_vgademo_on_fpga.magic.gds
string GDS_START 1096236
<< end >>

