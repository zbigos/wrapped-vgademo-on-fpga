* NGSPICE file created from wrapped_vgademo_on_fpga.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_8 abstract view
.subckt sky130_fd_sc_hd__ebufn_8 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_2 abstract view
.subckt sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_2 abstract view
.subckt sky130_fd_sc_hd__o32ai_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_4 abstract view
.subckt sky130_fd_sc_hd__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_1 abstract view
.subckt sky130_fd_sc_hd__o311ai_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

.subckt wrapped_vgademo_on_fpga active io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21]
+ io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29]
+ io_in[2] io_in[30] io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37]
+ io_in[3] io_in[4] io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10]
+ io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18]
+ io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25]
+ io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32]
+ io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5]
+ io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12]
+ io_out[13] io_out[14] io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1]
+ io_out[20] io_out[21] io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27]
+ io_out[28] io_out[29] io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34]
+ io_out[35] io_out[36] io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ io_out[8] io_out[9] la1_data_in[0] la1_data_in[10] la1_data_in[11] la1_data_in[12]
+ la1_data_in[13] la1_data_in[14] la1_data_in[15] la1_data_in[16] la1_data_in[17]
+ la1_data_in[18] la1_data_in[19] la1_data_in[1] la1_data_in[20] la1_data_in[21] la1_data_in[22]
+ la1_data_in[23] la1_data_in[24] la1_data_in[25] la1_data_in[26] la1_data_in[27]
+ la1_data_in[28] la1_data_in[29] la1_data_in[2] la1_data_in[30] la1_data_in[31] la1_data_in[3]
+ la1_data_in[4] la1_data_in[5] la1_data_in[6] la1_data_in[7] la1_data_in[8] la1_data_in[9]
+ la1_data_out[0] la1_data_out[10] la1_data_out[11] la1_data_out[12] la1_data_out[13]
+ la1_data_out[14] la1_data_out[15] la1_data_out[16] la1_data_out[17] la1_data_out[18]
+ la1_data_out[19] la1_data_out[1] la1_data_out[20] la1_data_out[21] la1_data_out[22]
+ la1_data_out[23] la1_data_out[24] la1_data_out[25] la1_data_out[26] la1_data_out[27]
+ la1_data_out[28] la1_data_out[29] la1_data_out[2] la1_data_out[30] la1_data_out[31]
+ la1_data_out[3] la1_data_out[4] la1_data_out[5] la1_data_out[6] la1_data_out[7]
+ la1_data_out[8] la1_data_out[9] la1_oenb[0] la1_oenb[10] la1_oenb[11] la1_oenb[12]
+ la1_oenb[13] la1_oenb[14] la1_oenb[15] la1_oenb[16] la1_oenb[17] la1_oenb[18] la1_oenb[19]
+ la1_oenb[1] la1_oenb[20] la1_oenb[21] la1_oenb[22] la1_oenb[23] la1_oenb[24] la1_oenb[25]
+ la1_oenb[26] la1_oenb[27] la1_oenb[28] la1_oenb[29] la1_oenb[2] la1_oenb[30] la1_oenb[31]
+ la1_oenb[3] la1_oenb[4] la1_oenb[5] la1_oenb[6] la1_oenb[7] la1_oenb[8] la1_oenb[9]
+ vccd1 vssd1 wb_clk_i
XFILLER_100_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7963_ _7963_/A vssd1 vssd1 vccd1 vccd1 _7963_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6914_ _6914_/A _6914_/B vssd1 vssd1 vccd1 vccd1 _6915_/B sky130_fd_sc_hd__and2_1
XFILLER_54_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7894_ _7893_/A _7893_/B _7893_/C vssd1 vssd1 vccd1 vccd1 _7946_/C sky130_fd_sc_hd__a21o_1
XFILLER_22_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6845_ _7099_/B _6845_/B vssd1 vssd1 vccd1 vccd1 _6845_/X sky130_fd_sc_hd__and2b_1
XFILLER_62_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6776_ _6784_/A vssd1 vssd1 vccd1 vccd1 _7443_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_22_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5727_ _5727_/A _5772_/B vssd1 vssd1 vccd1 vccd1 _5756_/A sky130_fd_sc_hd__xnor2_1
X_8515_ _8515_/A _8515_/B _8515_/C _8515_/D vssd1 vssd1 vccd1 vccd1 _8515_/X sky130_fd_sc_hd__and4_1
X_8446_ _7771_/A _7771_/C _7871_/X vssd1 vssd1 vccd1 vccd1 _8448_/A sky130_fd_sc_hd__a21o_1
X_5658_ _6028_/B vssd1 vssd1 vccd1 vccd1 _6193_/A sky130_fd_sc_hd__clkbuf_2
X_4609_ _8588_/Q _4610_/C _4608_/Y vssd1 vssd1 vccd1 vccd1 _8588_/D sky130_fd_sc_hd__a21oi_1
X_8377_ _8377_/A _8377_/B vssd1 vssd1 vccd1 vccd1 _8378_/B sky130_fd_sc_hd__xor2_1
X_5589_ _8658_/Q _6570_/B vssd1 vssd1 vccd1 vccd1 _5589_/X sky130_fd_sc_hd__and2b_1
X_7328_ _7328_/A _7328_/B vssd1 vssd1 vccd1 vccd1 _7439_/A sky130_fd_sc_hd__xnor2_1
XFILLER_89_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7259_ _7259_/A _7259_/B vssd1 vssd1 vccd1 vccd1 _7260_/B sky130_fd_sc_hd__nand2_1
XFILLER_58_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4960_ _4960_/A _4960_/B vssd1 vssd1 vccd1 vccd1 _4960_/X sky130_fd_sc_hd__or2_1
X_4891_ _4891_/A _4990_/A _4891_/C vssd1 vssd1 vccd1 vccd1 _4950_/B sky130_fd_sc_hd__or3_1
XFILLER_44_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6630_ _8701_/Q _8618_/Q vssd1 vssd1 vccd1 vccd1 _6659_/B sky130_fd_sc_hd__or2b_1
XFILLER_20_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6561_ _7060_/A vssd1 vssd1 vccd1 vccd1 _7335_/A sky130_fd_sc_hd__buf_2
X_8300_ _8239_/A _8300_/B vssd1 vssd1 vccd1 vccd1 _8300_/X sky130_fd_sc_hd__and2b_1
X_5512_ _5892_/A vssd1 vssd1 vccd1 vccd1 _5788_/A sky130_fd_sc_hd__inv_2
X_6492_ _8697_/Q vssd1 vssd1 vccd1 vccd1 _6536_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_8_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8231_ _8231_/A _8415_/B vssd1 vssd1 vccd1 vccd1 _8232_/B sky130_fd_sc_hd__nand2_1
X_5443_ _5874_/A vssd1 vssd1 vccd1 vccd1 _6020_/A sky130_fd_sc_hd__clkbuf_2
X_8162_ _8256_/B _8162_/B vssd1 vssd1 vccd1 vccd1 _8163_/B sky130_fd_sc_hd__nor2_2
X_5374_ _5374_/A _5374_/B _5389_/A vssd1 vssd1 vccd1 vccd1 _5374_/X sky130_fd_sc_hd__or3b_1
X_7113_ _7113_/A _7113_/B vssd1 vssd1 vccd1 vccd1 _7113_/Y sky130_fd_sc_hd__nor2_1
XFILLER_86_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8093_ _8094_/A _8094_/B vssd1 vssd1 vccd1 vccd1 _8186_/A sky130_fd_sc_hd__or2_1
XFILLER_101_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7044_ _6948_/X _6949_/Y _7042_/X _7043_/Y vssd1 vssd1 vccd1 vccd1 _7299_/A sky130_fd_sc_hd__o211a_1
XFILLER_86_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7946_ _7946_/A _7946_/B _7946_/C vssd1 vssd1 vccd1 vccd1 _7946_/X sky130_fd_sc_hd__and3_1
X_7877_ _7775_/A _7768_/B _7775_/B _7876_/X _7728_/A vssd1 vssd1 vccd1 vccd1 _7888_/A
+ sky130_fd_sc_hd__o311a_1
X_6828_ _6848_/A _6848_/B vssd1 vssd1 vccd1 vccd1 _6839_/B sky130_fd_sc_hd__and2_1
XFILLER_50_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6759_ _6759_/A _7324_/A vssd1 vssd1 vccd1 vccd1 _6804_/C sky130_fd_sc_hd__xnor2_2
XFILLER_12_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8429_ _8429_/A _8429_/B vssd1 vssd1 vccd1 vccd1 _8497_/B sky130_fd_sc_hd__xor2_1
XFILLER_2_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8745__12 vssd1 vssd1 vccd1 vccd1 _8745__12/HI _8840_/A sky130_fd_sc_hd__conb_1
XFILLER_53_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5090_ _5062_/C _5085_/X _5109_/D _5089_/X vssd1 vssd1 vccd1 vccd1 _5090_/X sky130_fd_sc_hd__o22a_1
XFILLER_78_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7800_ _8724_/Q _7906_/B vssd1 vssd1 vccd1 vccd1 _8051_/A sky130_fd_sc_hd__or2b_1
X_5992_ _5992_/A _5992_/B vssd1 vssd1 vccd1 vccd1 _6001_/A sky130_fd_sc_hd__nor2_2
XFILLER_91_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4943_ _4964_/B vssd1 vssd1 vccd1 vccd1 _5192_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_52_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7731_ _8206_/A _7839_/A _7796_/C _8122_/B vssd1 vssd1 vccd1 vccd1 _7841_/B sky130_fd_sc_hd__o211ai_2
X_7662_ _7662_/A _7661_/X vssd1 vssd1 vccd1 vccd1 _7725_/A sky130_fd_sc_hd__or2b_1
X_6613_ _6730_/A _6730_/B _7332_/A vssd1 vssd1 vccd1 vccd1 _6744_/A sky130_fd_sc_hd__a21o_1
X_4874_ _4877_/B vssd1 vssd1 vccd1 vccd1 _5196_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_20_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7593_ _7592_/Y _7590_/A _8543_/S vssd1 vssd1 vccd1 vccd1 _7594_/B sky130_fd_sc_hd__mux2_1
X_6544_ _7537_/C _6543_/C _6639_/A vssd1 vssd1 vccd1 vccd1 _6545_/C sky130_fd_sc_hd__o21ai_1
X_6475_ _8715_/Q _6500_/A _7532_/B vssd1 vssd1 vccd1 vccd1 _6475_/X sky130_fd_sc_hd__a21o_1
X_5426_ _5426_/A _5426_/B vssd1 vssd1 vccd1 vccd1 _5432_/B sky130_fd_sc_hd__or2_1
X_8214_ _8137_/A _8211_/B _8136_/B _8213_/Y vssd1 vssd1 vccd1 vccd1 _8237_/A sky130_fd_sc_hd__o31ai_4
XFILLER_99_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5357_ _8652_/Q _5358_/B vssd1 vssd1 vccd1 vccd1 _5359_/B sky130_fd_sc_hd__or2_1
X_8145_ _8145_/A vssd1 vssd1 vccd1 vccd1 _8150_/A sky130_fd_sc_hd__inv_2
X_5288_ _8638_/Q vssd1 vssd1 vccd1 vccd1 _6466_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_8076_ _8076_/A _8076_/B _8076_/C vssd1 vssd1 vccd1 vccd1 _8077_/B sky130_fd_sc_hd__nor3_1
XINSDIODE2_4 _4464_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7027_ _7027_/A _7027_/B vssd1 vssd1 vccd1 vccd1 _7036_/A sky130_fd_sc_hd__nand2_1
XFILLER_74_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7929_ _7928_/A _7928_/B _7928_/C vssd1 vssd1 vccd1 vccd1 _7929_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_43_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4590_ _8582_/Q _8581_/Q _8583_/Q vssd1 vssd1 vccd1 vccd1 _4591_/C sky130_fd_sc_hd__a21o_1
X_6260_ _6260_/A _6260_/B vssd1 vssd1 vccd1 vccd1 _6261_/B sky130_fd_sc_hd__xnor2_1
X_5211_ _5153_/A _5208_/X _5210_/X vssd1 vssd1 vccd1 vccd1 _5211_/X sky130_fd_sc_hd__o21a_1
X_6191_ _6191_/A _6191_/B vssd1 vssd1 vccd1 vccd1 _6191_/Y sky130_fd_sc_hd__nand2_1
X_5142_ _5207_/B _5229_/B _5109_/D _5173_/A vssd1 vssd1 vccd1 vccd1 _5143_/C sky130_fd_sc_hd__o31a_1
XFILLER_96_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5073_ _5073_/A _5078_/C _5072_/X vssd1 vssd1 vccd1 vccd1 _5073_/X sky130_fd_sc_hd__or3b_1
XFILLER_84_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8901_ _8901_/A _4461_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[0] sky130_fd_sc_hd__ebufn_8
XFILLER_92_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8832_ _8832_/A _4334_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[1] sky130_fd_sc_hd__ebufn_8
XFILLER_80_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5975_ _6168_/A _6238_/B _5974_/Y vssd1 vssd1 vccd1 vccd1 _5976_/B sky130_fd_sc_hd__a21oi_2
XFILLER_40_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8694_ _8695_/CLK _8694_/D vssd1 vssd1 vccd1 vccd1 _8694_/Q sky130_fd_sc_hd__dfxtp_1
X_4926_ _4942_/A _4979_/A vssd1 vssd1 vccd1 vccd1 _4927_/D sky130_fd_sc_hd__or2_1
XFILLER_33_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7714_ _7773_/A _8130_/A vssd1 vssd1 vccd1 vccd1 _8122_/B sky130_fd_sc_hd__nand2_2
X_4857_ _5127_/A _5233_/C vssd1 vssd1 vccd1 vccd1 _5120_/B sky130_fd_sc_hd__or2_1
X_7645_ _7645_/A _7644_/X vssd1 vssd1 vccd1 vccd1 _7656_/B sky130_fd_sc_hd__nor2b_2
XFILLER_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7576_ _7652_/A _7617_/B vssd1 vssd1 vccd1 vccd1 _7613_/A sky130_fd_sc_hd__nand2_1
X_6527_ _6522_/B _6524_/B _6520_/Y vssd1 vssd1 vccd1 vccd1 _6528_/C sky130_fd_sc_hd__a21oi_2
X_4788_ _4787_/A _5263_/B _4752_/X _4787_/Y vssd1 vssd1 vccd1 vccd1 _4789_/B sky130_fd_sc_hd__o2bb2a_1
X_6458_ _6458_/A vssd1 vssd1 vccd1 vccd1 _8692_/D sky130_fd_sc_hd__clkbuf_1
X_6389_ _8693_/Q _6388_/X _8694_/Q vssd1 vssd1 vccd1 vccd1 _6390_/B sky130_fd_sc_hd__a21o_1
X_5409_ _5404_/B _5397_/X _5398_/X _5408_/Y vssd1 vssd1 vccd1 vccd1 _8659_/D sky130_fd_sc_hd__a22o_1
XFILLER_87_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8128_ _8203_/A _8203_/B vssd1 vssd1 vccd1 vccd1 _8133_/A sky130_fd_sc_hd__nand2_1
XFILLER_102_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8059_ _8514_/A _8474_/A _8059_/C vssd1 vssd1 vccd1 vccd1 _8060_/A sky130_fd_sc_hd__or3_1
XFILLER_28_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5760_ _6028_/B vssd1 vssd1 vccd1 vccd1 _5944_/A sky130_fd_sc_hd__inv_2
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4711_ _4711_/A _4711_/B vssd1 vssd1 vccd1 vccd1 _4711_/X sky130_fd_sc_hd__or2_1
X_5691_ _5754_/B _5691_/B vssd1 vssd1 vccd1 vccd1 _5850_/A sky130_fd_sc_hd__nand2_1
X_7430_ _7430_/A _7430_/B vssd1 vssd1 vccd1 vccd1 _7432_/C sky130_fd_sc_hd__and2_1
X_4642_ _8599_/Q _4643_/C _4641_/Y vssd1 vssd1 vccd1 vccd1 _8599_/D sky130_fd_sc_hd__a21oi_1
XFILLER_30_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7361_ _7361_/A _6964_/B vssd1 vssd1 vccd1 vccd1 _7362_/C sky130_fd_sc_hd__or2b_1
X_4573_ _8592_/Q _8591_/Q _8594_/Q _8593_/Q vssd1 vssd1 vccd1 vccd1 _4577_/A sky130_fd_sc_hd__or4_1
X_7292_ _7293_/A _7292_/B vssd1 vssd1 vccd1 vccd1 _7295_/C sky130_fd_sc_hd__nand2_1
X_6312_ _6312_/A _6312_/B vssd1 vssd1 vccd1 vccd1 _6312_/X sky130_fd_sc_hd__xor2_1
X_6243_ _5493_/A _5493_/C _5491_/B vssd1 vssd1 vccd1 vccd1 _6245_/A sky130_fd_sc_hd__a21oi_1
XFILLER_69_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6174_ _6174_/A _6174_/B vssd1 vssd1 vccd1 vccd1 _6270_/B sky130_fd_sc_hd__xnor2_1
X_5125_ _4692_/A _5104_/X _5110_/X _5124_/X _4711_/B vssd1 vssd1 vccd1 vccd1 _5125_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_69_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5056_ _5056_/A _5056_/B vssd1 vssd1 vccd1 vccd1 _5056_/Y sky130_fd_sc_hd__nand2_1
XFILLER_84_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5958_ _5958_/A _5958_/B vssd1 vssd1 vccd1 vccd1 _5960_/C sky130_fd_sc_hd__xnor2_1
X_4909_ _4993_/A _5202_/C vssd1 vssd1 vccd1 vccd1 _5220_/B sky130_fd_sc_hd__or2_2
XFILLER_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8677_ _8677_/CLK _8677_/D vssd1 vssd1 vccd1 vccd1 _8677_/Q sky130_fd_sc_hd__dfxtp_1
X_5889_ _5889_/A _5889_/B vssd1 vssd1 vccd1 vccd1 _5983_/B sky130_fd_sc_hd__xnor2_1
XFILLER_21_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7628_ _8615_/Q _8718_/Q vssd1 vssd1 vccd1 vccd1 _7629_/A sky130_fd_sc_hd__or2b_1
X_7559_ _8716_/Q vssd1 vssd1 vccd1 vccd1 _8560_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6930_ _6932_/A _6854_/B _6929_/Y vssd1 vssd1 vccd1 vccd1 _7027_/A sky130_fd_sc_hd__o21bai_1
XFILLER_54_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6861_ _7039_/A _6861_/B vssd1 vssd1 vccd1 vccd1 _6862_/B sky130_fd_sc_hd__or2_1
XFILLER_81_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6792_ _6792_/A _6792_/B vssd1 vssd1 vccd1 vccd1 _6792_/Y sky130_fd_sc_hd__nand2_1
XFILLER_62_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8600_ _8600_/CLK _8600_/D vssd1 vssd1 vccd1 vccd1 _8600_/Q sky130_fd_sc_hd__dfxtp_1
X_5812_ _5812_/A vssd1 vssd1 vccd1 vccd1 _5970_/B sky130_fd_sc_hd__buf_2
XFILLER_62_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5743_ _5837_/B _6174_/A vssd1 vssd1 vccd1 vccd1 _5743_/Y sky130_fd_sc_hd__nand2_1
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8531_ _8531_/A _8727_/Q vssd1 vssd1 vccd1 vccd1 _8531_/Y sky130_fd_sc_hd__nor2_1
X_8462_ _8462_/A _8462_/B vssd1 vssd1 vccd1 vccd1 _8463_/B sky130_fd_sc_hd__xnor2_1
X_5674_ _6028_/A _5967_/A _5673_/Y vssd1 vssd1 vccd1 vccd1 _6033_/A sky130_fd_sc_hd__or3b_1
X_7413_ _7443_/B _7413_/B vssd1 vssd1 vccd1 vccd1 _7414_/S sky130_fd_sc_hd__nand2_1
X_4625_ _4628_/C _4625_/B vssd1 vssd1 vccd1 vccd1 _8593_/D sky130_fd_sc_hd__nor2_1
X_8393_ _8393_/A _8393_/B vssd1 vssd1 vccd1 vccd1 _8394_/B sky130_fd_sc_hd__nor2_1
X_7344_ _7344_/A vssd1 vssd1 vccd1 vccd1 _7345_/B sky130_fd_sc_hd__inv_2
X_4556_ _4556_/A vssd1 vssd1 vccd1 vccd1 _8885_/A sky130_fd_sc_hd__clkbuf_1
X_7275_ _7275_/A _7276_/B vssd1 vssd1 vccd1 vccd1 _7279_/B sky130_fd_sc_hd__xnor2_1
X_4487_ _4845_/B vssd1 vssd1 vccd1 vccd1 _4848_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6226_ _6226_/A _6226_/B vssd1 vssd1 vccd1 vccd1 _6227_/B sky130_fd_sc_hd__and2_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6157_ _6157_/A vssd1 vssd1 vccd1 vccd1 _6303_/A sky130_fd_sc_hd__inv_2
X_5108_ _5222_/B _5202_/D vssd1 vssd1 vccd1 vccd1 _5109_/C sky130_fd_sc_hd__or2_2
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6088_ _6148_/A _6148_/B _6087_/Y vssd1 vssd1 vccd1 vccd1 _6152_/A sky130_fd_sc_hd__o21a_1
X_5039_ _5218_/A _5096_/C vssd1 vssd1 vccd1 vccd1 _5043_/A sky130_fd_sc_hd__or2_1
XFILLER_72_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8729_ _8735_/CLK _8729_/D vssd1 vssd1 vccd1 vccd1 _8729_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8790__57 vssd1 vssd1 vccd1 vccd1 _8790__57/HI _8899_/A sky130_fd_sc_hd__conb_1
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4410_ _4413_/A vssd1 vssd1 vccd1 vccd1 _4410_/Y sky130_fd_sc_hd__inv_2
X_5390_ _5425_/B _5386_/X _5389_/Y _5279_/X vssd1 vssd1 vccd1 vccd1 _8656_/D sky130_fd_sc_hd__o211a_1
XFILLER_99_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4341_ _4344_/A vssd1 vssd1 vccd1 vccd1 _4341_/Y sky130_fd_sc_hd__inv_2
X_7060_ _7060_/A _7060_/B vssd1 vssd1 vccd1 vccd1 _7067_/A sky130_fd_sc_hd__or2_1
X_6011_ _6011_/A _6011_/B vssd1 vssd1 vccd1 vccd1 _6012_/B sky130_fd_sc_hd__xnor2_1
XFILLER_39_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7962_ _8119_/A vssd1 vssd1 vccd1 vccd1 _8044_/A sky130_fd_sc_hd__buf_2
X_6913_ _6914_/A _6914_/B vssd1 vssd1 vccd1 vccd1 _7033_/A sky130_fd_sc_hd__nor2_1
XFILLER_54_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7893_ _7893_/A _7893_/B _7893_/C vssd1 vssd1 vccd1 vccd1 _7946_/B sky130_fd_sc_hd__nand3_1
XFILLER_23_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6844_ _7095_/A _7095_/B vssd1 vssd1 vccd1 vccd1 _7096_/A sky130_fd_sc_hd__nand2_1
XFILLER_22_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6775_ _6775_/A _6892_/A vssd1 vssd1 vccd1 vccd1 _6784_/A sky130_fd_sc_hd__xnor2_1
XFILLER_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5726_ _5726_/A _5726_/B vssd1 vssd1 vccd1 vccd1 _5772_/B sky130_fd_sc_hd__xor2_2
XFILLER_22_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8514_ _8514_/A _8514_/B vssd1 vssd1 vccd1 vccd1 _8514_/X sky130_fd_sc_hd__or2_1
X_8445_ _8407_/A _8407_/B _8405_/A vssd1 vssd1 vccd1 vccd1 _8453_/A sky130_fd_sc_hd__o21a_1
X_5657_ _5728_/A _5728_/B vssd1 vssd1 vccd1 vccd1 _5669_/A sky130_fd_sc_hd__xnor2_1
X_4608_ _8588_/Q _4610_/C _4607_/X vssd1 vssd1 vccd1 vccd1 _4608_/Y sky130_fd_sc_hd__o21ai_1
X_8376_ _8292_/A _8292_/B _8375_/X vssd1 vssd1 vccd1 vccd1 _8377_/B sky130_fd_sc_hd__a21oi_1
X_5588_ _8658_/Q _6570_/B vssd1 vssd1 vccd1 vccd1 _5638_/B sky130_fd_sc_hd__xnor2_4
X_7327_ _7327_/A _7436_/B vssd1 vssd1 vccd1 vccd1 _7328_/B sky130_fd_sc_hd__xor2_1
X_4539_ _4781_/A _4864_/A _4808_/A _4765_/A vssd1 vssd1 vccd1 vccd1 _4660_/B sky130_fd_sc_hd__or4_1
XFILLER_104_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7258_ _7258_/A _7258_/B vssd1 vssd1 vccd1 vccd1 _7259_/B sky130_fd_sc_hd__nand2_1
XFILLER_77_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6209_ _6209_/A _6209_/B vssd1 vssd1 vccd1 vccd1 _6239_/B sky130_fd_sc_hd__xnor2_1
X_7189_ _7190_/A _7190_/B _7190_/C vssd1 vssd1 vccd1 vccd1 _7189_/Y sky130_fd_sc_hd__o21ai_1
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4890_ _4990_/A _4890_/B vssd1 vssd1 vccd1 vccd1 _5233_/B sky130_fd_sc_hd__nor2_2
XFILLER_32_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6560_ _6835_/A vssd1 vssd1 vccd1 vccd1 _7060_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5511_ _6019_/A _6019_/B _5510_/X vssd1 vssd1 vccd1 vccd1 _5552_/A sky130_fd_sc_hd__a21o_1
X_6491_ _6515_/A _6509_/A _6521_/A vssd1 vssd1 vccd1 vccd1 _6491_/Y sky130_fd_sc_hd__o21ai_1
X_8230_ _8231_/A _8415_/B vssd1 vssd1 vccd1 vccd1 _8341_/B sky130_fd_sc_hd__or2_1
X_5442_ _5474_/A vssd1 vssd1 vccd1 vccd1 _5874_/A sky130_fd_sc_hd__buf_2
X_8161_ _8161_/A _8161_/B vssd1 vssd1 vccd1 vccd1 _8162_/B sky130_fd_sc_hd__nor2_1
X_5373_ _5456_/A _6341_/A _8671_/Q vssd1 vssd1 vccd1 vccd1 _5374_/B sky130_fd_sc_hd__o21a_1
XFILLER_99_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7112_ _7112_/A _7112_/B vssd1 vssd1 vccd1 vccd1 _7156_/B sky130_fd_sc_hd__xnor2_1
X_8092_ _8180_/A _8092_/B vssd1 vssd1 vccd1 vccd1 _8094_/B sky130_fd_sc_hd__nand2_1
X_7043_ _7302_/A _7042_/B _7042_/C vssd1 vssd1 vccd1 vccd1 _7043_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_86_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7945_ _7945_/A _7945_/B _7945_/C vssd1 vssd1 vccd1 vccd1 _7945_/X sky130_fd_sc_hd__and3_1
X_7876_ _7876_/A _6596_/B vssd1 vssd1 vccd1 vccd1 _7876_/X sky130_fd_sc_hd__or2b_1
X_6827_ _6826_/A _6826_/B _6826_/C vssd1 vssd1 vccd1 vccd1 _6848_/B sky130_fd_sc_hd__a21o_2
XFILLER_23_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6758_ _7000_/A vssd1 vssd1 vccd1 vccd1 _7324_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_7_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6689_ _6689_/A vssd1 vssd1 vccd1 vccd1 _6689_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5709_ _5709_/A _5777_/B vssd1 vssd1 vccd1 vccd1 _5716_/A sky130_fd_sc_hd__xnor2_1
X_8428_ _8491_/A _8428_/B vssd1 vssd1 vccd1 vccd1 _8429_/B sky130_fd_sc_hd__nor2_1
X_8359_ _8350_/A _8359_/B vssd1 vssd1 vccd1 vccd1 _8359_/X sky130_fd_sc_hd__and2b_1
XFILLER_104_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8760__27 vssd1 vssd1 vccd1 vccd1 _8760__27/HI _8855_/A sky130_fd_sc_hd__conb_1
XFILLER_41_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_12_0_wb_clk_i clkbuf_3_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8714_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5991_ _5872_/B _5993_/A _6001_/B _5569_/X vssd1 vssd1 vccd1 vccd1 _6202_/A sky130_fd_sc_hd__a31o_1
X_4942_ _4942_/A vssd1 vssd1 vccd1 vccd1 _5215_/A sky130_fd_sc_hd__buf_2
XFILLER_64_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7730_ _8321_/A _7887_/A vssd1 vssd1 vccd1 vccd1 _7839_/A sky130_fd_sc_hd__nor2_1
X_7661_ _7661_/A _7835_/B _7661_/C vssd1 vssd1 vccd1 vccd1 _7661_/X sky130_fd_sc_hd__or3_1
X_6612_ _7146_/A vssd1 vssd1 vccd1 vccd1 _7465_/A sky130_fd_sc_hd__clkbuf_4
X_4873_ _4876_/A _4906_/A _4872_/X vssd1 vssd1 vccd1 vccd1 _4877_/B sky130_fd_sc_hd__o21ai_1
XFILLER_60_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7592_ _8718_/Q _7592_/B vssd1 vssd1 vccd1 vccd1 _7592_/Y sky130_fd_sc_hd__xnor2_1
X_6543_ _6639_/A _7548_/B _6543_/C vssd1 vssd1 vccd1 vccd1 _6545_/B sky130_fd_sc_hd__or3_1
X_6474_ _7526_/B vssd1 vssd1 vccd1 vccd1 _7532_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_8213_ _8213_/A _8213_/B vssd1 vssd1 vccd1 vccd1 _8213_/Y sky130_fd_sc_hd__nand2_1
X_5425_ _5426_/A _5425_/B vssd1 vssd1 vccd1 vccd1 _5427_/C sky130_fd_sc_hd__nand2_1
X_5356_ _5358_/B _5356_/B vssd1 vssd1 vccd1 vccd1 _8651_/D sky130_fd_sc_hd__nor2_1
X_8144_ _8192_/A _8192_/B vssd1 vssd1 vccd1 vccd1 _8163_/A sky130_fd_sc_hd__xor2_2
XFILLER_101_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5287_ _8635_/Q _8634_/Q vssd1 vssd1 vccd1 vccd1 _5301_/A sky130_fd_sc_hd__or2_1
XFILLER_87_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8075_ _8076_/A _8076_/C _8076_/B vssd1 vssd1 vccd1 vccd1 _8161_/A sky130_fd_sc_hd__o21a_1
XINSDIODE2_5 _8574_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7026_ _6920_/A _6920_/B _7025_/X vssd1 vssd1 vccd1 vccd1 _7300_/B sky130_fd_sc_hd__a21o_1
XFILLER_101_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7928_ _7928_/A _7928_/B _7928_/C vssd1 vssd1 vccd1 vccd1 _7928_/X sky130_fd_sc_hd__and3_1
XFILLER_43_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7859_ _8118_/A _7859_/B _7859_/C vssd1 vssd1 vccd1 vccd1 _7950_/B sky130_fd_sc_hd__and3_1
XFILLER_11_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8805__72 vssd1 vssd1 vccd1 vccd1 _8805__72/HI _8914_/A sky130_fd_sc_hd__conb_1
XFILLER_65_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5210_ _5227_/D _5210_/B _5210_/C vssd1 vssd1 vccd1 vccd1 _5210_/X sky130_fd_sc_hd__or3_1
X_6190_ _6255_/A _6190_/B vssd1 vssd1 vccd1 vccd1 _6198_/A sky130_fd_sc_hd__nor2_2
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5141_ _5137_/X _5139_/X _5140_/X vssd1 vssd1 vccd1 vccd1 _5141_/X sky130_fd_sc_hd__o21a_1
XFILLER_96_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5072_ _4522_/A _5068_/Y _5069_/X _5070_/Y _5248_/A vssd1 vssd1 vccd1 vccd1 _5072_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_69_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8900_ _8900_/A _4427_/Y vssd1 vssd1 vccd1 vccd1 io_out[37] sky130_fd_sc_hd__ebufn_8
XFILLER_64_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8831_ _8831_/A _4464_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[0] sky130_fd_sc_hd__ebufn_8
XFILLER_25_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5974_ _6194_/A _5974_/B vssd1 vssd1 vccd1 vccd1 _5974_/Y sky130_fd_sc_hd__nor2_1
X_7713_ _7713_/A _7713_/B vssd1 vssd1 vccd1 vccd1 _8130_/A sky130_fd_sc_hd__xnor2_4
X_8693_ _8695_/CLK _8693_/D vssd1 vssd1 vccd1 vccd1 _8693_/Q sky130_fd_sc_hd__dfxtp_1
X_4925_ _4914_/A _5136_/B _4924_/X vssd1 vssd1 vccd1 vccd1 _4927_/C sky130_fd_sc_hd__o21a_1
X_4856_ _5138_/A _5114_/A vssd1 vssd1 vccd1 vccd1 _5233_/C sky130_fd_sc_hd__or2_2
XFILLER_60_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7644_ _7644_/A _8618_/Q vssd1 vssd1 vccd1 vccd1 _7644_/X sky130_fd_sc_hd__or2_1
X_7575_ _8722_/Q vssd1 vssd1 vccd1 vccd1 _7652_/A sky130_fd_sc_hd__inv_2
X_6526_ _6531_/A _6526_/B vssd1 vssd1 vccd1 vccd1 _6534_/A sky130_fd_sc_hd__nand2_1
X_4787_ _4787_/A _4787_/B vssd1 vssd1 vccd1 vccd1 _4787_/Y sky130_fd_sc_hd__xnor2_1
X_6457_ _6459_/B _6457_/B _6457_/C vssd1 vssd1 vccd1 vccd1 _6458_/A sky130_fd_sc_hd__and3b_1
X_6388_ _8690_/Q _6455_/B _6395_/A _6387_/X _8692_/Q vssd1 vssd1 vccd1 vccd1 _6388_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5408_ _5408_/A _5408_/B vssd1 vssd1 vccd1 vccd1 _5408_/Y sky130_fd_sc_hd__xnor2_1
X_5339_ _6468_/C _8644_/Q _5332_/B _8646_/Q vssd1 vssd1 vccd1 vccd1 _5340_/C sky130_fd_sc_hd__a31o_1
X_8127_ _8213_/A _8213_/B vssd1 vssd1 vccd1 vccd1 _8137_/A sky130_fd_sc_hd__xnor2_2
XFILLER_102_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8058_ _8052_/A _7836_/C _8054_/A vssd1 vssd1 vccd1 vccd1 _8059_/C sky130_fd_sc_hd__a21oi_1
X_7009_ _7060_/A _7009_/B vssd1 vssd1 vccd1 vccd1 _7010_/B sky130_fd_sc_hd__or2_1
XFILLER_47_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4710_ _4710_/A vssd1 vssd1 vccd1 vccd1 _4711_/B sky130_fd_sc_hd__clkbuf_2
X_5690_ _5754_/B _5691_/B _5690_/C vssd1 vssd1 vccd1 vccd1 _5769_/A sky130_fd_sc_hd__and3_1
X_4641_ _8599_/Q _4643_/C _4612_/B vssd1 vssd1 vccd1 vccd1 _4641_/Y sky130_fd_sc_hd__o21ai_1
X_7360_ _7356_/A _7447_/B _7359_/C vssd1 vssd1 vccd1 vccd1 _7362_/B sky130_fd_sc_hd__a21o_1
X_4572_ _8584_/Q _8583_/Q _8586_/Q _8585_/Q vssd1 vssd1 vccd1 vccd1 _4578_/B sky130_fd_sc_hd__or4_1
X_7291_ _7291_/A _7163_/B vssd1 vssd1 vccd1 vccd1 _7295_/B sky130_fd_sc_hd__or2b_1
X_6311_ _6311_/A _6311_/B vssd1 vssd1 vccd1 vccd1 _6311_/Y sky130_fd_sc_hd__nand2_1
XFILLER_89_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6242_ _6242_/A _6242_/B vssd1 vssd1 vccd1 vccd1 _6250_/A sky130_fd_sc_hd__xor2_1
X_6173_ _6172_/Y _5969_/B _5967_/X vssd1 vssd1 vccd1 vccd1 _6175_/A sky130_fd_sc_hd__a21boi_1
X_5124_ _5017_/C _5123_/X _5065_/A vssd1 vssd1 vccd1 vccd1 _5124_/X sky130_fd_sc_hd__o21a_1
XFILLER_84_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5055_ _4697_/X _5052_/X _5054_/X vssd1 vssd1 vccd1 vccd1 _5056_/B sky130_fd_sc_hd__o21ai_1
XFILLER_84_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8796__63 vssd1 vssd1 vccd1 vccd1 _8796__63/HI _8905_/A sky130_fd_sc_hd__conb_1
XFILLER_65_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5957_ _5957_/A _6179_/B vssd1 vssd1 vccd1 vccd1 _5958_/B sky130_fd_sc_hd__xnor2_1
XFILLER_13_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8676_ _8677_/CLK _8676_/D vssd1 vssd1 vccd1 vccd1 _8676_/Q sky130_fd_sc_hd__dfxtp_1
X_4908_ _5046_/A _5018_/A vssd1 vssd1 vccd1 vccd1 _5202_/C sky130_fd_sc_hd__or2_2
XFILLER_80_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5888_ _5896_/A _6218_/B vssd1 vssd1 vccd1 vccd1 _5889_/B sky130_fd_sc_hd__xnor2_1
X_7627_ _7577_/X _7625_/Y _7626_/Y vssd1 vssd1 vccd1 vccd1 _8724_/D sky130_fd_sc_hd__a21oi_1
X_4839_ _4839_/A _4839_/B _4848_/C _4848_/A vssd1 vssd1 vccd1 vccd1 _4990_/B sky130_fd_sc_hd__or4b_4
X_7558_ _8732_/Q vssd1 vssd1 vccd1 vccd1 _8553_/A sky130_fd_sc_hd__inv_2
X_6509_ _6509_/A _6536_/B vssd1 vssd1 vccd1 vccd1 _6511_/B sky130_fd_sc_hd__xor2_1
X_7489_ _7487_/X _7488_/Y _7489_/S vssd1 vssd1 vccd1 vccd1 _7489_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6860_ _7039_/A _6861_/B vssd1 vssd1 vccd1 vccd1 _6862_/A sky130_fd_sc_hd__nand2_1
X_6791_ _6792_/A _6792_/B vssd1 vssd1 vccd1 vccd1 _6791_/X sky130_fd_sc_hd__or2_1
X_5811_ _5811_/A _5948_/B vssd1 vssd1 vccd1 vccd1 _5812_/A sky130_fd_sc_hd__and2_1
X_5742_ _5742_/A _6030_/B vssd1 vssd1 vccd1 vccd1 _5837_/B sky130_fd_sc_hd__nand2_1
XFILLER_22_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8530_ _8533_/B _8529_/Y _8525_/A _8525_/B vssd1 vssd1 vccd1 vccd1 _8530_/X sky130_fd_sc_hd__a211o_1
X_5673_ _5673_/A _5673_/B vssd1 vssd1 vccd1 vccd1 _5673_/Y sky130_fd_sc_hd__xnor2_1
X_8461_ _8461_/A _8461_/B vssd1 vssd1 vccd1 vccd1 _8462_/B sky130_fd_sc_hd__or2_1
X_7412_ _7412_/A _7412_/B vssd1 vssd1 vccd1 vccd1 _7418_/A sky130_fd_sc_hd__xnor2_1
X_4624_ _8593_/Q _4623_/B _4607_/X vssd1 vssd1 vccd1 vccd1 _4625_/B sky130_fd_sc_hd__o21ai_1
X_8392_ _8392_/A _8392_/B _8392_/C vssd1 vssd1 vccd1 vccd1 _8393_/B sky130_fd_sc_hd__and3_1
X_7343_ _7341_/Y _7015_/B _7342_/Y vssd1 vssd1 vccd1 vccd1 _7344_/A sky130_fd_sc_hd__a21oi_1
X_4555_ _8631_/Q _4563_/B vssd1 vssd1 vccd1 vccd1 _4556_/A sky130_fd_sc_hd__and2_1
XFILLER_89_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7274_ _7274_/A _7274_/B vssd1 vssd1 vccd1 vccd1 _7276_/B sky130_fd_sc_hd__xor2_1
X_4486_ _8614_/Q vssd1 vssd1 vccd1 vccd1 _4845_/B sky130_fd_sc_hd__clkbuf_2
X_6225_ _6226_/A _6226_/B vssd1 vssd1 vccd1 vccd1 _6227_/A sky130_fd_sc_hd__nor2_1
XFILLER_97_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6156_ _6311_/A _6311_/B _6153_/X _6155_/X vssd1 vssd1 vccd1 vccd1 _6306_/B sky130_fd_sc_hd__a31o_1
XFILLER_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5107_ _5107_/A _5188_/B _5107_/C vssd1 vssd1 vccd1 vccd1 _5202_/D sky130_fd_sc_hd__or3_2
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6087_ _6087_/A _6087_/B vssd1 vssd1 vccd1 vccd1 _6087_/Y sky130_fd_sc_hd__nand2_1
X_5038_ _5038_/A _5248_/B vssd1 vssd1 vccd1 vccd1 _5096_/C sky130_fd_sc_hd__or2_2
XFILLER_72_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6989_ _6989_/A _6989_/B _6989_/C vssd1 vssd1 vccd1 vccd1 _7347_/C sky130_fd_sc_hd__and3_1
XFILLER_53_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8728_ _8735_/CLK _8728_/D vssd1 vssd1 vccd1 vccd1 _8728_/Q sky130_fd_sc_hd__dfxtp_1
X_8659_ _8732_/CLK _8659_/D vssd1 vssd1 vccd1 vccd1 _8659_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4340_ _4344_/A vssd1 vssd1 vccd1 vccd1 _4340_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6010_ _6010_/A _6165_/B vssd1 vssd1 vccd1 vccd1 _6011_/B sky130_fd_sc_hd__xnor2_1
XFILLER_67_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7961_ _8515_/C _8130_/B vssd1 vssd1 vccd1 vccd1 _8119_/A sky130_fd_sc_hd__or2_1
X_8766__33 vssd1 vssd1 vccd1 vccd1 _8766__33/HI _8861_/A sky130_fd_sc_hd__conb_1
X_6912_ _6995_/A _6995_/B vssd1 vssd1 vccd1 vccd1 _6918_/A sky130_fd_sc_hd__xnor2_1
X_7892_ _7980_/A _7892_/B vssd1 vssd1 vccd1 vccd1 _7893_/C sky130_fd_sc_hd__and2b_1
X_6843_ _7409_/B _6833_/Y _6842_/Y vssd1 vssd1 vccd1 vccd1 _7095_/B sky130_fd_sc_hd__o21ai_1
XFILLER_62_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6774_ _7169_/B _6773_/X _6774_/S vssd1 vssd1 vccd1 vccd1 _6892_/A sky130_fd_sc_hd__mux2_2
XFILLER_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5725_ _5987_/A _5722_/X _5824_/A vssd1 vssd1 vccd1 vccd1 _5726_/B sky130_fd_sc_hd__a21oi_1
X_8513_ _8514_/A _8514_/B vssd1 vssd1 vccd1 vccd1 _8518_/A sky130_fd_sc_hd__nand2_1
X_5656_ _5729_/A _5729_/B vssd1 vssd1 vccd1 vccd1 _5728_/B sky130_fd_sc_hd__xor2_1
X_8444_ _8418_/A _8418_/B _8443_/Y vssd1 vssd1 vccd1 vccd1 _8454_/A sky130_fd_sc_hd__a21oi_1
X_4607_ _4607_/A vssd1 vssd1 vccd1 vccd1 _4607_/X sky130_fd_sc_hd__clkbuf_2
X_8375_ _8293_/B _8375_/B vssd1 vssd1 vccd1 vccd1 _8375_/X sky130_fd_sc_hd__and2b_1
X_5587_ _5587_/A vssd1 vssd1 vccd1 vccd1 _5642_/A sky130_fd_sc_hd__clkbuf_4
X_7326_ _7427_/A _7326_/B vssd1 vssd1 vccd1 vccd1 _7436_/B sky130_fd_sc_hd__nand2_1
XFILLER_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4538_ _4900_/A _4957_/A _4749_/A vssd1 vssd1 vccd1 vccd1 _4754_/B sky130_fd_sc_hd__a21o_1
X_4469_ _6553_/B vssd1 vssd1 vccd1 vccd1 _4480_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_7257_ _7274_/A _7274_/B _7256_/A vssd1 vssd1 vccd1 vccd1 _7260_/A sky130_fd_sc_hd__a21oi_2
XFILLER_104_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6208_ _6253_/A _6253_/B _6207_/X vssd1 vssd1 vccd1 vccd1 _6209_/B sky130_fd_sc_hd__o21ba_1
X_7188_ _7188_/A _7188_/B _7188_/C vssd1 vssd1 vccd1 vccd1 _7188_/Y sky130_fd_sc_hd__nor3_2
XFILLER_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6139_ _6295_/A _6298_/A vssd1 vssd1 vccd1 vccd1 _6299_/B sky130_fd_sc_hd__or2_1
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5510_ _6071_/A _5872_/A _5510_/C vssd1 vssd1 vccd1 vccd1 _5510_/X sky130_fd_sc_hd__and3_1
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6490_ _8701_/Q vssd1 vssd1 vccd1 vccd1 _6521_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5441_ _5540_/A _6316_/A vssd1 vssd1 vccd1 vccd1 _5474_/A sky130_fd_sc_hd__xor2_1
XFILLER_99_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8160_ _8161_/A _8161_/B vssd1 vssd1 vccd1 vccd1 _8256_/B sky130_fd_sc_hd__and2_1
X_5372_ _5456_/A _6341_/A _8668_/Q _6354_/A vssd1 vssd1 vccd1 vccd1 _5372_/X sky130_fd_sc_hd__a31o_1
X_7111_ _7151_/A _7151_/B vssd1 vssd1 vccd1 vccd1 _7112_/A sky130_fd_sc_hd__nand2_1
X_8091_ _8091_/A _8091_/B vssd1 vssd1 vccd1 vccd1 _8092_/B sky130_fd_sc_hd__or2_1
X_7042_ _7302_/A _7042_/B _7042_/C vssd1 vssd1 vccd1 vccd1 _7042_/X sky130_fd_sc_hd__or3_1
XFILLER_101_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7944_ _7846_/Y _8529_/A _7943_/X vssd1 vssd1 vccd1 vccd1 _8525_/A sky130_fd_sc_hd__a21oi_1
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7875_ _7875_/A _8204_/A vssd1 vssd1 vccd1 vccd1 _7963_/A sky130_fd_sc_hd__nor2_1
X_6826_ _6826_/A _6826_/B _6826_/C vssd1 vssd1 vccd1 vccd1 _6848_/A sky130_fd_sc_hd__nand3_4
XFILLER_11_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6757_ _6724_/A _6694_/B _6804_/A vssd1 vssd1 vccd1 vccd1 _6803_/B sky130_fd_sc_hd__a21bo_1
XFILLER_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5708_ _5708_/A _5795_/A vssd1 vssd1 vccd1 vccd1 _5777_/B sky130_fd_sc_hd__xor2_2
X_6688_ _6688_/A vssd1 vssd1 vccd1 vccd1 _6688_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_8427_ _8427_/A _8427_/B _8427_/C vssd1 vssd1 vccd1 vccd1 _8428_/B sky130_fd_sc_hd__nor3_1
X_5639_ _5652_/A vssd1 vssd1 vccd1 vccd1 _5859_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8358_ _8299_/A _8299_/B _8357_/X vssd1 vssd1 vccd1 vccd1 _8425_/A sky130_fd_sc_hd__a21oi_1
XFILLER_104_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7309_ _7196_/C _7007_/B _6916_/B vssd1 vssd1 vccd1 vccd1 _7312_/A sky130_fd_sc_hd__o21ai_2
X_8289_ _8289_/A _8289_/B vssd1 vssd1 vccd1 vccd1 _8362_/B sky130_fd_sc_hd__xnor2_1
XFILLER_104_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5990_ _5903_/A _5901_/X _5902_/A vssd1 vssd1 vccd1 vccd1 _6006_/A sky130_fd_sc_hd__a21o_1
XFILLER_91_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4941_ _5171_/C _5044_/C _4987_/B _4941_/D vssd1 vssd1 vccd1 vccd1 _4941_/X sky130_fd_sc_hd__or4_1
XFILLER_52_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4872_ _4903_/B _4879_/B _4917_/A vssd1 vssd1 vccd1 vccd1 _4872_/X sky130_fd_sc_hd__o21a_1
XFILLER_17_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7660_ _7813_/A _8281_/B _7661_/C vssd1 vssd1 vccd1 vccd1 _7662_/A sky130_fd_sc_hd__o21a_1
X_6611_ _7102_/A vssd1 vssd1 vccd1 vccd1 _7146_/A sky130_fd_sc_hd__buf_2
XFILLER_20_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7591_ _7591_/A _7591_/B vssd1 vssd1 vccd1 vccd1 _7592_/B sky130_fd_sc_hd__nand2_1
X_6542_ _6531_/A _6528_/C _6537_/B _6541_/X vssd1 vssd1 vccd1 vccd1 _6543_/C sky130_fd_sc_hd__o31a_1
X_6473_ _8696_/Q vssd1 vssd1 vccd1 vccd1 _7526_/B sky130_fd_sc_hd__inv_2
XFILLER_9_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8212_ _8316_/A _8212_/B vssd1 vssd1 vccd1 vccd1 _8238_/A sky130_fd_sc_hd__and2_1
X_5424_ _5398_/A _5422_/X _5433_/S _5397_/X _5432_/A vssd1 vssd1 vccd1 vccd1 _8661_/D
+ sky130_fd_sc_hd__a32o_1
X_8143_ _8143_/A _8143_/B vssd1 vssd1 vccd1 vccd1 _8192_/B sky130_fd_sc_hd__xnor2_2
XFILLER_99_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5355_ _8651_/Q _5354_/B _5311_/X vssd1 vssd1 vccd1 vccd1 _5356_/B sky130_fd_sc_hd__o21ai_1
XFILLER_101_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_6 _4545_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5286_ _8708_/Q _5271_/A _5285_/X _5279_/X vssd1 vssd1 vccd1 vccd1 _8633_/D sky130_fd_sc_hd__o211a_1
X_8074_ _8172_/A _8074_/B vssd1 vssd1 vccd1 vccd1 _8076_/B sky130_fd_sc_hd__and2b_1
X_7025_ _6919_/A _7025_/B vssd1 vssd1 vccd1 vccd1 _7025_/X sky130_fd_sc_hd__and2b_1
XFILLER_87_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7927_ _8020_/A _7927_/B vssd1 vssd1 vccd1 vccd1 _7928_/C sky130_fd_sc_hd__nor2_1
XFILLER_70_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7858_ _7780_/A _7780_/B _7857_/X vssd1 vssd1 vccd1 vccd1 _7883_/A sky130_fd_sc_hd__a21o_1
XFILLER_90_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6809_ _6745_/A _6747_/A _6745_/B _6602_/Y vssd1 vssd1 vccd1 vccd1 _6812_/A sky130_fd_sc_hd__a31o_1
XFILLER_23_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7789_ _7861_/A vssd1 vssd1 vccd1 vccd1 _8331_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8820__87 vssd1 vssd1 vccd1 vccd1 _8820__87/HI _8929_/A sky130_fd_sc_hd__conb_1
XFILLER_64_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5140_ _5120_/D _5118_/Y _5128_/X _4665_/A vssd1 vssd1 vccd1 vccd1 _5140_/X sky130_fd_sc_hd__o22a_1
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5071_ _5226_/A vssd1 vssd1 vccd1 vccd1 _5248_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_65_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5973_ _5973_/A _6174_/B vssd1 vssd1 vccd1 vccd1 _6238_/B sky130_fd_sc_hd__xnor2_2
XFILLER_25_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4924_ _4900_/A _4900_/B _4820_/X _4923_/X vssd1 vssd1 vccd1 vccd1 _4924_/X sky130_fd_sc_hd__a31o_1
XFILLER_52_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7712_ _7712_/A _7712_/B vssd1 vssd1 vccd1 vccd1 _7773_/A sky130_fd_sc_hd__xnor2_2
X_8692_ _8695_/CLK _8692_/D vssd1 vssd1 vccd1 vccd1 _8692_/Q sky130_fd_sc_hd__dfxtp_1
X_4855_ _5186_/C _5002_/B vssd1 vssd1 vccd1 vccd1 _5114_/A sky130_fd_sc_hd__or2_1
X_7643_ _7644_/A _7643_/B vssd1 vssd1 vccd1 vccd1 _7645_/A sky130_fd_sc_hd__and2_1
X_4786_ _4786_/A _4786_/B _4786_/C vssd1 vssd1 vccd1 vccd1 _4787_/B sky130_fd_sc_hd__and3_1
X_7574_ _7597_/A _7574_/B vssd1 vssd1 vccd1 vccd1 _7574_/Y sky130_fd_sc_hd__nand2_1
X_6525_ _6521_/A _5362_/X _6508_/X _6524_/Y vssd1 vssd1 vccd1 vccd1 _8701_/D sky130_fd_sc_hd__a22o_1
X_6456_ _8690_/Q _6455_/B _6450_/B _8692_/Q vssd1 vssd1 vccd1 vccd1 _6457_/C sky130_fd_sc_hd__a31o_1
XFILLER_69_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6387_ _8687_/Q _6385_/X _6446_/B vssd1 vssd1 vccd1 vccd1 _6387_/X sky130_fd_sc_hd__a21o_1
X_5407_ _5615_/A _5402_/B _5401_/A vssd1 vssd1 vccd1 vccd1 _5408_/B sky130_fd_sc_hd__o21a_1
XFILLER_102_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5338_ _8646_/Q _6468_/C _5338_/C vssd1 vssd1 vccd1 vccd1 _5345_/C sky130_fd_sc_hd__and3_1
X_8126_ _8126_/A _8126_/B vssd1 vssd1 vccd1 vccd1 _8213_/B sky130_fd_sc_hd__xnor2_1
X_8057_ _8057_/A vssd1 vssd1 vccd1 vccd1 _8474_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7008_ _7028_/A _6800_/A _7310_/A vssd1 vssd1 vccd1 vccd1 _7416_/A sky130_fd_sc_hd__mux2_1
XFILLER_75_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5269_ _8626_/Q _5276_/B vssd1 vssd1 vccd1 vccd1 _5269_/X sky130_fd_sc_hd__or2_1
XFILLER_47_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4640_ _4640_/A vssd1 vssd1 vccd1 vccd1 _8598_/D sky130_fd_sc_hd__clkbuf_1
X_6310_ _6311_/A _6311_/B vssd1 vssd1 vccd1 vccd1 _6310_/X sky130_fd_sc_hd__or2_1
X_4571_ _8582_/Q _8581_/Q vssd1 vssd1 vccd1 vccd1 _4587_/A sky130_fd_sc_hd__or2_1
X_7290_ _7481_/A _7481_/B _7479_/A _7478_/A vssd1 vssd1 vccd1 vccd1 _7475_/C sky130_fd_sc_hd__o211ai_2
X_6241_ _6221_/A _6215_/A _6221_/X _6223_/A vssd1 vssd1 vccd1 vccd1 _6242_/B sky130_fd_sc_hd__o22a_1
XFILLER_103_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6172_ _6172_/A vssd1 vssd1 vccd1 vccd1 _6172_/Y sky130_fd_sc_hd__inv_2
X_5123_ _5233_/C _5062_/C _5113_/X _5122_/X vssd1 vssd1 vccd1 vccd1 _5123_/X sky130_fd_sc_hd__o31a_1
XFILLER_69_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5054_ _5054_/A _5155_/B _5065_/D _5096_/C vssd1 vssd1 vccd1 vccd1 _5054_/X sky130_fd_sc_hd__or4_1
XFILLER_57_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5956_ _6193_/B _5956_/B vssd1 vssd1 vccd1 vccd1 _6179_/B sky130_fd_sc_hd__xnor2_1
XFILLER_40_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8675_ _8677_/CLK _8675_/D vssd1 vssd1 vccd1 vccd1 _8675_/Q sky130_fd_sc_hd__dfxtp_1
X_4907_ _4932_/A _5207_/D vssd1 vssd1 vccd1 vccd1 _5018_/A sky130_fd_sc_hd__or2_1
XFILLER_21_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5887_ _6218_/A _5794_/B _5782_/B _5872_/B vssd1 vssd1 vccd1 vccd1 _5983_/A sky130_fd_sc_hd__a22o_1
XFILLER_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4838_ _4955_/A _4956_/A vssd1 vssd1 vccd1 vccd1 _5054_/A sky130_fd_sc_hd__or2_2
X_7626_ _7577_/X _7625_/Y _4771_/X vssd1 vssd1 vccd1 vccd1 _7626_/Y sky130_fd_sc_hd__o21ai_1
X_4769_ _4769_/A vssd1 vssd1 vccd1 vccd1 _8616_/D sky130_fd_sc_hd__clkbuf_1
X_7557_ _8731_/Q _8540_/A _8732_/Q vssd1 vssd1 vccd1 vccd1 _7557_/X sky130_fd_sc_hd__o21a_1
X_6508_ _6508_/A vssd1 vssd1 vccd1 vccd1 _6508_/X sky130_fd_sc_hd__buf_2
X_7488_ _7488_/A vssd1 vssd1 vccd1 vccd1 _7488_/Y sky130_fd_sc_hd__clkinv_2
X_6439_ _6441_/B _6439_/B _6457_/B vssd1 vssd1 vccd1 vccd1 _6440_/A sky130_fd_sc_hd__and3b_1
XFILLER_20_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8109_ _8096_/A _8096_/B _8108_/X vssd1 vssd1 vccd1 vccd1 _8187_/A sky130_fd_sc_hd__a21oi_1
XFILLER_102_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6790_ _6790_/A _6790_/B vssd1 vssd1 vccd1 vccd1 _6819_/A sky130_fd_sc_hd__nor2_1
XFILLER_62_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5810_ _5810_/A vssd1 vssd1 vccd1 vccd1 _5827_/A sky130_fd_sc_hd__inv_2
XFILLER_22_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5741_ _5971_/A vssd1 vssd1 vccd1 vccd1 _6193_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8460_ _8460_/A _8460_/B vssd1 vssd1 vccd1 vccd1 _8462_/A sky130_fd_sc_hd__nor2_1
X_7411_ _7444_/A _7411_/B vssd1 vssd1 vccd1 vccd1 _7412_/B sky130_fd_sc_hd__xnor2_1
X_5672_ _5952_/A _6028_/B vssd1 vssd1 vccd1 vccd1 _5673_/B sky130_fd_sc_hd__nor2_1
X_4623_ _8593_/Q _4623_/B vssd1 vssd1 vccd1 vccd1 _4628_/C sky130_fd_sc_hd__and2_1
X_8391_ _8392_/A _8392_/B _8392_/C vssd1 vssd1 vccd1 vccd1 _8393_/A sky130_fd_sc_hd__a21oi_1
X_7342_ _7342_/A _7342_/B vssd1 vssd1 vccd1 vccd1 _7342_/Y sky130_fd_sc_hd__nor2_1
X_4554_ _4567_/B vssd1 vssd1 vccd1 vccd1 _4563_/B sky130_fd_sc_hd__clkbuf_1
X_7273_ _7283_/A _7273_/B vssd1 vssd1 vccd1 vccd1 _7278_/A sky130_fd_sc_hd__nand2_1
XFILLER_103_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4485_ _5634_/B vssd1 vssd1 vccd1 vccd1 _4787_/A sky130_fd_sc_hd__clkbuf_2
X_6224_ _6224_/A _6224_/B vssd1 vssd1 vccd1 vccd1 _6226_/B sky130_fd_sc_hd__xnor2_1
XFILLER_103_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6155_ _6307_/A _6154_/X _6307_/B vssd1 vssd1 vccd1 vccd1 _6155_/X sky130_fd_sc_hd__o21ba_1
X_5106_ _5215_/B _5106_/B _5106_/C _5229_/C vssd1 vssd1 vccd1 vccd1 _5106_/X sky130_fd_sc_hd__or4_1
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6086_ _6087_/A _6087_/B vssd1 vssd1 vccd1 vccd1 _6148_/B sky130_fd_sc_hd__xnor2_1
XFILLER_85_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5037_ _5037_/A _5233_/C vssd1 vssd1 vccd1 vccd1 _5248_/B sky130_fd_sc_hd__or2_1
XFILLER_38_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6988_ _7003_/A _6889_/B _6987_/X vssd1 vssd1 vccd1 vccd1 _6989_/C sky130_fd_sc_hd__a21o_1
XFILLER_80_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8727_ _8735_/CLK _8727_/D vssd1 vssd1 vccd1 vccd1 _8727_/Q sky130_fd_sc_hd__dfxtp_1
X_5939_ _5831_/X _5910_/B _5913_/B _5938_/X vssd1 vssd1 vccd1 vccd1 _5958_/A sky130_fd_sc_hd__a31o_1
XFILLER_40_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8658_ _8732_/CLK _8658_/D vssd1 vssd1 vccd1 vccd1 _8658_/Q sky130_fd_sc_hd__dfxtp_2
X_8589_ _8600_/CLK _8589_/D vssd1 vssd1 vccd1 vccd1 _8589_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7609_ _8721_/Q vssd1 vssd1 vccd1 vccd1 _7644_/A sky130_fd_sc_hd__inv_2
XFILLER_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7960_ _8217_/A _7960_/B vssd1 vssd1 vccd1 vccd1 _7965_/A sky130_fd_sc_hd__nand2_1
X_6911_ _6911_/A _6911_/B vssd1 vssd1 vccd1 vccd1 _6995_/B sky130_fd_sc_hd__xnor2_1
XFILLER_82_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7891_ _7891_/A _7891_/B _7891_/C vssd1 vssd1 vccd1 vccd1 _7892_/B sky130_fd_sc_hd__or3_1
X_6842_ _7072_/A _7072_/B vssd1 vssd1 vccd1 vccd1 _6842_/Y sky130_fd_sc_hd__nand2_1
XFILLER_90_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8781__48 vssd1 vssd1 vccd1 vccd1 _8781__48/HI _8890_/A sky130_fd_sc_hd__conb_1
X_6773_ _6625_/X _6688_/X _6689_/X _6670_/B _6876_/A vssd1 vssd1 vccd1 vccd1 _6773_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_22_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5724_ _5722_/X _5723_/X _5987_/A vssd1 vssd1 vccd1 vccd1 _5824_/A sky130_fd_sc_hd__a21oi_2
X_8512_ _8512_/A _8512_/B _8512_/C _8512_/D vssd1 vssd1 vccd1 vccd1 _8525_/B sky130_fd_sc_hd__or4_4
X_5655_ _5833_/A _6182_/A vssd1 vssd1 vccd1 vccd1 _5729_/B sky130_fd_sc_hd__xnor2_2
X_8443_ _8443_/A _8443_/B vssd1 vssd1 vccd1 vccd1 _8443_/Y sky130_fd_sc_hd__nor2_1
X_4606_ _4610_/C _4606_/B vssd1 vssd1 vccd1 vccd1 _8587_/D sky130_fd_sc_hd__nor2_1
X_8374_ _8374_/A _8374_/B vssd1 vssd1 vccd1 vccd1 _8377_/A sky130_fd_sc_hd__xnor2_1
X_7325_ _7369_/B _7324_/A vssd1 vssd1 vccd1 vccd1 _7326_/B sky130_fd_sc_hd__or2b_1
X_5586_ _8615_/Q _8657_/Q vssd1 vssd1 vccd1 vccd1 _5587_/A sky130_fd_sc_hd__or2b_1
X_4537_ _4834_/C vssd1 vssd1 vccd1 vccd1 _4957_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_104_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4468_ _8606_/Q vssd1 vssd1 vccd1 vccd1 _6553_/B sky130_fd_sc_hd__buf_2
X_7256_ _7256_/A _7256_/B vssd1 vssd1 vccd1 vccd1 _7274_/B sky130_fd_sc_hd__nor2_1
X_7187_ _7187_/A _7187_/B vssd1 vssd1 vccd1 vccd1 _7188_/C sky130_fd_sc_hd__xnor2_1
X_6207_ _6253_/A _6204_/Y _6206_/X vssd1 vssd1 vccd1 vccd1 _6207_/X sky130_fd_sc_hd__o21a_1
X_4399_ _4400_/A vssd1 vssd1 vccd1 vccd1 _4399_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_58_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6138_ _6297_/A _6322_/A vssd1 vssd1 vccd1 vccd1 _6298_/A sky130_fd_sc_hd__nand2_1
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6069_ _6069_/A _6069_/B vssd1 vssd1 vccd1 vccd1 _6073_/A sky130_fd_sc_hd__xor2_1
XFILLER_26_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5440_ _8669_/Q _8606_/Q vssd1 vssd1 vccd1 vccd1 _6316_/A sky130_fd_sc_hd__xnor2_4
XFILLER_8_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5371_ _6353_/A _6353_/B vssd1 vssd1 vccd1 vccd1 _6354_/A sky130_fd_sc_hd__nand2_1
XFILLER_99_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7110_ _7113_/A _7113_/B vssd1 vssd1 vccd1 vccd1 _7156_/A sky130_fd_sc_hd__xor2_1
X_8090_ _8091_/A _8091_/B vssd1 vssd1 vccd1 vccd1 _8180_/A sky130_fd_sc_hd__nand2_2
XFILLER_99_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7041_ _7041_/A _7041_/B vssd1 vssd1 vccd1 vccd1 _7042_/C sky130_fd_sc_hd__xnor2_1
X_8826__93 vssd1 vssd1 vccd1 vccd1 _8826__93/HI _8935_/A sky130_fd_sc_hd__conb_1
XFILLER_79_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7943_ _8102_/B _7943_/B vssd1 vssd1 vccd1 vccd1 _7943_/X sky130_fd_sc_hd__xor2_1
XFILLER_70_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7874_ _8130_/B vssd1 vssd1 vccd1 vccd1 _8204_/A sky130_fd_sc_hd__clkbuf_2
X_6825_ _6825_/A _6825_/B vssd1 vssd1 vccd1 vccd1 _6826_/C sky130_fd_sc_hd__nand2_1
Xclkbuf_3_7_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
X_6756_ _6856_/A _6756_/B vssd1 vssd1 vccd1 vccd1 _6763_/A sky130_fd_sc_hd__and2_1
XFILLER_50_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5707_ _5873_/A _5884_/B vssd1 vssd1 vccd1 vccd1 _5795_/A sky130_fd_sc_hd__nor2_2
X_6687_ _6734_/A vssd1 vssd1 vccd1 vccd1 _7254_/A sky130_fd_sc_hd__clkbuf_2
X_8426_ _8427_/A _8427_/B _8427_/C vssd1 vssd1 vccd1 vccd1 _8491_/A sky130_fd_sc_hd__o21a_1
X_5638_ _5642_/A _5638_/B vssd1 vssd1 vccd1 vccd1 _5652_/A sky130_fd_sc_hd__xor2_2
XFILLER_88_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8357_ _8298_/A _8357_/B vssd1 vssd1 vccd1 vccd1 _8357_/X sky130_fd_sc_hd__and2b_1
X_5569_ _5569_/A vssd1 vssd1 vccd1 vccd1 _5569_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7308_ _7034_/A _7033_/B _7033_/A vssd1 vssd1 vccd1 vccd1 _7316_/A sky130_fd_sc_hd__a21oi_1
XFILLER_88_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8288_ _8365_/B _8288_/B vssd1 vssd1 vccd1 vccd1 _8289_/B sky130_fd_sc_hd__nand2_1
X_7239_ _7430_/A _6841_/A _7065_/X vssd1 vssd1 vccd1 vccd1 _7239_/X sky130_fd_sc_hd__o21a_1
XFILLER_77_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4940_ _4923_/X _5115_/A _4939_/X vssd1 vssd1 vccd1 vccd1 _4941_/D sky130_fd_sc_hd__o21a_1
X_4871_ _4876_/A _4920_/B _4830_/A _4903_/B _4870_/Y vssd1 vssd1 vccd1 vccd1 _4917_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_60_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8751__18 vssd1 vssd1 vccd1 vccd1 _8751__18/HI _8846_/A sky130_fd_sc_hd__conb_1
X_6610_ _6914_/A vssd1 vssd1 vccd1 vccd1 _7102_/A sky130_fd_sc_hd__buf_2
XFILLER_60_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7590_ _7590_/A _8717_/Q vssd1 vssd1 vccd1 vccd1 _7591_/B sky130_fd_sc_hd__or2b_1
X_6541_ _6541_/A _6541_/B vssd1 vssd1 vccd1 vccd1 _6541_/X sky130_fd_sc_hd__or2_1
X_6472_ _8637_/Q _8636_/Q _6472_/C _6472_/D vssd1 vssd1 vccd1 vccd1 _6500_/A sky130_fd_sc_hd__and4_2
X_8211_ _8211_/A _8211_/B _8211_/C vssd1 vssd1 vccd1 vccd1 _8212_/B sky130_fd_sc_hd__or3_1
X_5423_ _5427_/A _5423_/B _5423_/C vssd1 vssd1 vccd1 vccd1 _5433_/S sky130_fd_sc_hd__nand3_1
X_5354_ _8651_/Q _5354_/B vssd1 vssd1 vccd1 vccd1 _5358_/B sky130_fd_sc_hd__and2_1
X_8142_ _8402_/A _8195_/B vssd1 vssd1 vccd1 vccd1 _8143_/B sky130_fd_sc_hd__xnor2_2
XINSDIODE2_7 _6503_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5285_ _8633_/Q _5285_/B vssd1 vssd1 vccd1 vccd1 _5285_/X sky130_fd_sc_hd__or2_1
XFILLER_59_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8073_ _8072_/A _8284_/A _8072_/D _8072_/C vssd1 vssd1 vccd1 vccd1 _8074_/B sky130_fd_sc_hd__a31o_1
XFILLER_101_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7024_ _7403_/A _6939_/B _7023_/X vssd1 vssd1 vccd1 vccd1 _7041_/A sky130_fd_sc_hd__a21o_1
XFILLER_95_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7926_ _7926_/A _7926_/B vssd1 vssd1 vccd1 vccd1 _7927_/B sky130_fd_sc_hd__and2_1
XFILLER_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7857_ _8208_/A _8217_/A _7857_/C vssd1 vssd1 vccd1 vccd1 _7857_/X sky130_fd_sc_hd__and3_1
X_6808_ _6797_/A _6914_/A _6916_/B vssd1 vssd1 vccd1 vccd1 _7007_/B sky130_fd_sc_hd__a21bo_1
X_7788_ _7955_/C _7955_/D vssd1 vssd1 vccd1 vccd1 _7861_/A sky130_fd_sc_hd__nor2_1
XFILLER_51_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6739_ _6914_/A _7000_/A vssd1 vssd1 vccd1 vccd1 _7127_/A sky130_fd_sc_hd__xor2_4
X_8409_ _8331_/A _8411_/S _8332_/B _8410_/B vssd1 vssd1 vccd1 vccd1 _8412_/A sky130_fd_sc_hd__a22o_1
XFILLER_74_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5070_ _5106_/B _5207_/D vssd1 vssd1 vccd1 vccd1 _5070_/Y sky130_fd_sc_hd__nor2_1
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5972_ _5974_/B _6194_/B vssd1 vssd1 vccd1 vccd1 _6174_/B sky130_fd_sc_hd__and2_1
X_4923_ _4923_/A vssd1 vssd1 vccd1 vccd1 _4923_/X sky130_fd_sc_hd__buf_2
X_7711_ _7711_/A _7711_/B vssd1 vssd1 vccd1 vccd1 _8139_/A sky130_fd_sc_hd__xnor2_4
X_8691_ _8695_/CLK _8691_/D vssd1 vssd1 vccd1 vccd1 _8691_/Q sky130_fd_sc_hd__dfxtp_1
X_4854_ _5007_/A _4963_/B vssd1 vssd1 vccd1 vccd1 _5002_/B sky130_fd_sc_hd__or2_1
XFILLER_60_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7642_ _7642_/A _7642_/B vssd1 vssd1 vccd1 vccd1 _7656_/A sky130_fd_sc_hd__nand2_2
X_4785_ _4785_/A vssd1 vssd1 vccd1 vccd1 _8558_/A sky130_fd_sc_hd__clkbuf_4
X_7573_ _7590_/A _8718_/Q _8721_/Q vssd1 vssd1 vccd1 vccd1 _7574_/B sky130_fd_sc_hd__a21oi_1
X_6524_ _6524_/A _6524_/B vssd1 vssd1 vccd1 vccd1 _6524_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_20_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6455_ _8692_/Q _6455_/B _6455_/C vssd1 vssd1 vccd1 vccd1 _6459_/B sky130_fd_sc_hd__and3_1
X_6386_ _8688_/Q vssd1 vssd1 vccd1 vccd1 _6446_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_5406_ _5406_/A _5406_/B vssd1 vssd1 vccd1 vccd1 _5408_/A sky130_fd_sc_hd__nor2_1
X_5337_ _6468_/C _5338_/C _5336_/Y vssd1 vssd1 vccd1 vccd1 _8645_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8125_ _8224_/A _8323_/A _8225_/A vssd1 vssd1 vccd1 vccd1 _8126_/B sky130_fd_sc_hd__o21a_1
X_5268_ _8667_/Q _5258_/X _5266_/X _5267_/X vssd1 vssd1 vccd1 vccd1 _8625_/D sky130_fd_sc_hd__o211a_1
X_8056_ _8085_/B _8087_/B vssd1 vssd1 vccd1 vccd1 _8061_/A sky130_fd_sc_hd__or2b_1
XFILLER_87_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7007_ _7054_/B _7007_/B vssd1 vssd1 vccd1 vccd1 _7013_/A sky130_fd_sc_hd__xnor2_1
X_5199_ _5199_/A _5200_/A _5199_/C _5229_/B vssd1 vssd1 vccd1 vccd1 _5199_/X sky130_fd_sc_hd__or4_1
XFILLER_56_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7909_ _7804_/A _7804_/B _7910_/A _7798_/B vssd1 vssd1 vccd1 vccd1 _8008_/A sky130_fd_sc_hd__o211a_1
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8889_ _8889_/A _4403_/Y vssd1 vssd1 vccd1 vccd1 io_out[26] sky130_fd_sc_hd__ebufn_8
XFILLER_24_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4570_ _7499_/A vssd1 vssd1 vccd1 vccd1 _8531_/A sky130_fd_sc_hd__clkbuf_2
X_6240_ _6213_/A _6213_/B _6239_/Y vssd1 vssd1 vccd1 vccd1 _6251_/A sky130_fd_sc_hd__o21a_1
X_6171_ _6171_/A _6171_/B vssd1 vssd1 vccd1 vccd1 _6176_/A sky130_fd_sc_hd__nand2_1
X_5122_ _4665_/A _5118_/Y _5120_/X _5230_/D vssd1 vssd1 vccd1 vccd1 _5122_/X sky130_fd_sc_hd__o22a_1
XFILLER_97_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5053_ _5053_/A _5166_/A vssd1 vssd1 vccd1 vccd1 _5065_/D sky130_fd_sc_hd__or2_1
XFILLER_65_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5955_ _5955_/A _5955_/B vssd1 vssd1 vccd1 vccd1 _5957_/A sky130_fd_sc_hd__xnor2_1
XFILLER_40_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4906_ _4906_/A _5047_/B vssd1 vssd1 vccd1 vccd1 _5207_/D sky130_fd_sc_hd__nor2_2
X_5886_ _6218_/B _5708_/A _5795_/A _5795_/B vssd1 vssd1 vccd1 vccd1 _5891_/A sky130_fd_sc_hd__a22o_1
X_8674_ _8674_/CLK _8674_/D vssd1 vssd1 vccd1 vccd1 _8674_/Q sky130_fd_sc_hd__dfxtp_1
X_4837_ _4891_/C _4837_/B vssd1 vssd1 vccd1 vccd1 _4956_/A sky130_fd_sc_hd__nor2_1
X_7625_ _8578_/A _7625_/B vssd1 vssd1 vccd1 vccd1 _7625_/Y sky130_fd_sc_hd__nor2_1
XFILLER_21_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4768_ _4779_/B _7550_/A _4768_/C vssd1 vssd1 vccd1 vccd1 _4769_/A sky130_fd_sc_hd__and3b_1
X_7556_ _8730_/Q vssd1 vssd1 vccd1 vccd1 _8540_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4699_ _5064_/A vssd1 vssd1 vccd1 vccd1 _5056_/A sky130_fd_sc_hd__clkbuf_2
X_6507_ _6507_/A vssd1 vssd1 vccd1 vccd1 _6508_/A sky130_fd_sc_hd__clkbuf_2
X_7487_ _7395_/X _7394_/X _7488_/A vssd1 vssd1 vccd1 vccd1 _7487_/X sky130_fd_sc_hd__a21o_1
X_6438_ _6437_/B _8684_/Q _6431_/A _8686_/Q vssd1 vssd1 vccd1 vccd1 _6439_/B sky130_fd_sc_hd__a31o_1
XFILLER_0_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8108_ _8083_/B _8108_/B vssd1 vssd1 vccd1 vccd1 _8108_/X sky130_fd_sc_hd__and2b_1
X_6369_ _6369_/A _6372_/B vssd1 vssd1 vccd1 vccd1 _6370_/B sky130_fd_sc_hd__or2_1
XFILLER_102_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8039_ _8116_/A _8039_/B vssd1 vssd1 vccd1 vccd1 _8040_/B sky130_fd_sc_hd__and2_1
XFILLER_48_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8787__54 vssd1 vssd1 vccd1 vccd1 _8787__54/HI _8896_/A sky130_fd_sc_hd__conb_1
XFILLER_16_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5740_ _5944_/B _6030_/B vssd1 vssd1 vccd1 vccd1 _5971_/A sky130_fd_sc_hd__nand2_1
XFILLER_22_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7410_ _7338_/A _7338_/B _7409_/Y _7337_/B vssd1 vssd1 vccd1 vccd1 _7411_/B sky130_fd_sc_hd__a22o_1
X_5671_ _5948_/A _5948_/B vssd1 vssd1 vccd1 vccd1 _5673_/A sky130_fd_sc_hd__nand2_1
XFILLER_30_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4622_ _4622_/A vssd1 vssd1 vccd1 vccd1 _8592_/D sky130_fd_sc_hd__clkbuf_1
X_8390_ _8390_/A _8460_/B vssd1 vssd1 vccd1 vccd1 _8392_/C sky130_fd_sc_hd__xnor2_1
X_7341_ _7342_/A _7342_/B vssd1 vssd1 vccd1 vccd1 _7341_/Y sky130_fd_sc_hd__nand2_1
X_4553_ _4553_/A vssd1 vssd1 vccd1 vccd1 _8884_/A sky130_fd_sc_hd__clkbuf_1
X_7272_ _7272_/A _7272_/B vssd1 vssd1 vccd1 vccd1 _7273_/B sky130_fd_sc_hd__or2_1
X_4484_ _7906_/B vssd1 vssd1 vccd1 vccd1 _5634_/B sky130_fd_sc_hd__clkbuf_2
X_6223_ _6223_/A _6223_/B vssd1 vssd1 vccd1 vccd1 _6224_/B sky130_fd_sc_hd__xnor2_1
XFILLER_97_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6154_ _6299_/A _6151_/A _6154_/C _6154_/D vssd1 vssd1 vccd1 vccd1 _6154_/X sky130_fd_sc_hd__and4bb_1
X_5105_ _5212_/A _5107_/C _5109_/B vssd1 vssd1 vccd1 vccd1 _5229_/C sky130_fd_sc_hd__or3_2
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6085_ _6085_/A _6085_/B vssd1 vssd1 vccd1 vccd1 _6087_/B sky130_fd_sc_hd__xor2_1
XFILLER_85_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5036_ _5097_/A vssd1 vssd1 vccd1 vccd1 _5218_/A sky130_fd_sc_hd__clkbuf_2
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6987_ _6897_/A _6987_/B vssd1 vssd1 vccd1 vccd1 _6987_/X sky130_fd_sc_hd__and2b_1
XFILLER_41_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5938_ _6238_/A _5938_/B vssd1 vssd1 vccd1 vccd1 _5938_/X sky130_fd_sc_hd__and2b_1
XFILLER_25_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8726_ _8735_/CLK _8726_/D vssd1 vssd1 vccd1 vccd1 _8726_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5869_ _5869_/A _5869_/B vssd1 vssd1 vccd1 vccd1 _5907_/A sky130_fd_sc_hd__xor2_2
X_8657_ _8674_/CLK _8657_/D vssd1 vssd1 vccd1 vccd1 _8657_/Q sky130_fd_sc_hd__dfxtp_1
X_8588_ _8600_/CLK _8588_/D vssd1 vssd1 vccd1 vccd1 _8588_/Q sky130_fd_sc_hd__dfxtp_1
X_7608_ _7652_/A _7618_/B vssd1 vssd1 vccd1 vccd1 _7613_/B sky130_fd_sc_hd__or2_1
X_7539_ _7540_/A _8696_/Q vssd1 vssd1 vccd1 vccd1 _7539_/Y sky130_fd_sc_hd__nand2_1
XFILLER_5_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_4_9_0_wb_clk_i clkbuf_4_9_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _8677_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_97_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6910_ _7004_/A _7327_/A vssd1 vssd1 vccd1 vccd1 _6911_/B sky130_fd_sc_hd__xor2_1
X_7890_ _7891_/A _7891_/B _7891_/C vssd1 vssd1 vccd1 vccd1 _7980_/A sky130_fd_sc_hd__o21a_1
XFILLER_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6841_ _6841_/A _6857_/A vssd1 vssd1 vccd1 vccd1 _7072_/B sky130_fd_sc_hd__and2_1
XFILLER_62_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6772_ _6980_/A _6774_/S _6708_/X vssd1 vssd1 vccd1 vccd1 _7364_/B sky130_fd_sc_hd__o21ai_4
XFILLER_50_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8511_ _8501_/X _8502_/Y _8505_/X _8508_/Y _8510_/Y vssd1 vssd1 vccd1 vccd1 _8512_/D
+ sky130_fd_sc_hd__a2111o_1
X_5723_ _5723_/A _5581_/B vssd1 vssd1 vccd1 vccd1 _5723_/X sky130_fd_sc_hd__or2b_1
X_5654_ _5737_/A vssd1 vssd1 vccd1 vccd1 _6182_/A sky130_fd_sc_hd__clkbuf_4
X_8442_ _8442_/A _8442_/B vssd1 vssd1 vccd1 vccd1 _8466_/A sky130_fd_sc_hd__xnor2_1
X_8373_ _8373_/A _8469_/B vssd1 vssd1 vccd1 vccd1 _8374_/B sky130_fd_sc_hd__xnor2_1
XFILLER_30_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4605_ _8587_/Q _4603_/A _4595_/X vssd1 vssd1 vccd1 vccd1 _4606_/B sky130_fd_sc_hd__o21ai_1
X_7324_ _7324_/A _7369_/B vssd1 vssd1 vccd1 vccd1 _7427_/A sky130_fd_sc_hd__or2b_1
X_5585_ _5694_/A _5694_/B vssd1 vssd1 vccd1 vccd1 _6047_/A sky130_fd_sc_hd__xor2_1
X_4536_ _8612_/Q vssd1 vssd1 vccd1 vccd1 _4834_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_104_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7255_ _7254_/A _7254_/B _7254_/C vssd1 vssd1 vccd1 vccd1 _7256_/B sky130_fd_sc_hd__a21oi_1
X_4467_ _7677_/B vssd1 vssd1 vccd1 vccd1 _6603_/B sky130_fd_sc_hd__buf_2
X_7186_ _7185_/A _7185_/C _7185_/B vssd1 vssd1 vccd1 vccd1 _7188_/B sky130_fd_sc_hd__a21oi_1
X_4398_ _4400_/A vssd1 vssd1 vccd1 vccd1 _4398_/Y sky130_fd_sc_hd__inv_2
X_6206_ _5892_/A _6020_/Y _5997_/A vssd1 vssd1 vccd1 vccd1 _6206_/X sky130_fd_sc_hd__a21o_1
X_6137_ _6321_/A _6321_/B vssd1 vssd1 vccd1 vccd1 _6322_/A sky130_fd_sc_hd__nor2_1
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6068_ _6075_/A _6075_/B _6082_/B vssd1 vssd1 vccd1 vccd1 _6148_/A sky130_fd_sc_hd__or3b_1
X_8757__24 vssd1 vssd1 vccd1 vccd1 _8757__24/HI _8852_/A sky130_fd_sc_hd__conb_1
X_5019_ _5171_/A _5227_/A vssd1 vssd1 vccd1 vccd1 _5062_/C sky130_fd_sc_hd__or2_2
XFILLER_73_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8709_ _8715_/CLK _8709_/D vssd1 vssd1 vccd1 vccd1 _8709_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5370_ _8671_/Q vssd1 vssd1 vccd1 vccd1 _6353_/A sky130_fd_sc_hd__inv_2
X_7040_ _7300_/B _7040_/B vssd1 vssd1 vccd1 vccd1 _7041_/B sky130_fd_sc_hd__xnor2_1
XFILLER_101_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7942_ _8101_/A _8102_/A vssd1 vssd1 vccd1 vccd1 _7943_/B sky130_fd_sc_hd__nand2_1
XFILLER_82_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7873_ _7952_/B vssd1 vssd1 vccd1 vccd1 _8130_/B sky130_fd_sc_hd__clkbuf_1
X_6824_ _8714_/Q _6598_/A vssd1 vssd1 vccd1 vccd1 _6825_/B sky130_fd_sc_hd__or2b_1
X_6755_ _6841_/A _7196_/C _7102_/A vssd1 vssd1 vccd1 vccd1 _6756_/B sky130_fd_sc_hd__o21ai_1
X_5706_ _5532_/A _5708_/A _5564_/B _5574_/A vssd1 vssd1 vccd1 vccd1 _5778_/A sky130_fd_sc_hd__a22oi_2
X_6686_ _6780_/A _6685_/C _6793_/C vssd1 vssd1 vccd1 vccd1 _6697_/B sky130_fd_sc_hd__a21o_1
X_8425_ _8425_/A _8425_/B vssd1 vssd1 vccd1 vccd1 _8427_/C sky130_fd_sc_hd__xor2_1
X_5637_ _5941_/A _5944_/B vssd1 vssd1 vccd1 vccd1 _5962_/A sky130_fd_sc_hd__nand2_2
X_8356_ _8353_/A _8356_/B vssd1 vssd1 vccd1 vccd1 _8427_/B sky130_fd_sc_hd__and2b_1
X_5568_ _6108_/A _5992_/B vssd1 vssd1 vccd1 vccd1 _5569_/A sky130_fd_sc_hd__nor2_1
X_7307_ _7017_/A _7017_/B _7306_/X vssd1 vssd1 vccd1 vccd1 _7406_/B sky130_fd_sc_hd__a21bo_1
X_4519_ _8602_/Q vssd1 vssd1 vccd1 vccd1 _5245_/A sky130_fd_sc_hd__clkbuf_2
X_8287_ _8365_/A _8069_/A _8365_/C vssd1 vssd1 vccd1 vccd1 _8288_/B sky130_fd_sc_hd__mux2_1
XFILLER_104_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7238_ _7238_/A _7238_/B vssd1 vssd1 vccd1 vccd1 _7258_/A sky130_fd_sc_hd__xnor2_1
X_5499_ _5499_/A _5539_/C vssd1 vssd1 vccd1 vccd1 _5500_/B sky130_fd_sc_hd__xnor2_1
XFILLER_77_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7169_ _7169_/A _7169_/B vssd1 vssd1 vccd1 vccd1 _7170_/B sky130_fd_sc_hd__nand2_1
XFILLER_58_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4870_ _5185_/B _5190_/B vssd1 vssd1 vccd1 vccd1 _4870_/Y sky130_fd_sc_hd__nor2_1
XFILLER_60_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6540_ _8704_/Q vssd1 vssd1 vccd1 vccd1 _6639_/A sky130_fd_sc_hd__inv_2
XFILLER_20_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6471_ _5301_/A _6471_/B _6471_/C _6471_/D vssd1 vssd1 vccd1 vccd1 _6472_/D sky130_fd_sc_hd__and4b_1
X_5422_ _5427_/A _5423_/B _5423_/C vssd1 vssd1 vccd1 vccd1 _5422_/X sky130_fd_sc_hd__a21o_1
X_8210_ _8211_/A _8211_/B _8211_/C vssd1 vssd1 vccd1 vccd1 _8316_/A sky130_fd_sc_hd__o21ai_4
X_5353_ _5354_/B _5353_/B vssd1 vssd1 vccd1 vccd1 _8650_/D sky130_fd_sc_hd__nor2_1
X_8141_ _8041_/A _8041_/B _8040_/A vssd1 vssd1 vccd1 vccd1 _8195_/B sky130_fd_sc_hd__a21o_1
XFILLER_87_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5284_ _8707_/Q _5271_/A _5283_/X _5279_/X vssd1 vssd1 vccd1 vccd1 _8632_/D sky130_fd_sc_hd__o211a_1
X_8072_ _8072_/A _8284_/A _8072_/C _8072_/D vssd1 vssd1 vccd1 vccd1 _8172_/A sky130_fd_sc_hd__and4_1
X_7023_ _6938_/B _7023_/B vssd1 vssd1 vccd1 vccd1 _7023_/X sky130_fd_sc_hd__and2b_1
XINSDIODE2_8 _4942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7925_ _7926_/A _7926_/B vssd1 vssd1 vccd1 vccd1 _8020_/A sky130_fd_sc_hd__nor2_1
XFILLER_63_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7856_ _7859_/C vssd1 vssd1 vccd1 vccd1 _8217_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_23_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6807_ _6807_/A _7443_/A vssd1 vssd1 vccd1 vccd1 _6916_/B sky130_fd_sc_hd__nand2_2
XFILLER_51_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4999_ _4999_/A _5236_/C vssd1 vssd1 vccd1 vccd1 _5067_/C sky130_fd_sc_hd__or2_1
XFILLER_11_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7787_ _7960_/B vssd1 vssd1 vccd1 vccd1 _8203_/B sky130_fd_sc_hd__clkbuf_2
X_6738_ _7370_/A _7076_/B vssd1 vssd1 vccd1 vccd1 _6742_/A sky130_fd_sc_hd__or2b_1
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6669_ _6669_/A vssd1 vssd1 vccd1 vccd1 _6694_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_8408_ _8343_/A _8343_/B _8342_/A vssd1 vssd1 vccd1 vccd1 _8418_/A sky130_fd_sc_hd__a21o_1
XFILLER_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8339_ _8415_/B _8415_/C vssd1 vssd1 vccd1 vccd1 _8413_/B sky130_fd_sc_hd__xnor2_1
XFILLER_2_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8737__4 vssd1 vssd1 vccd1 vccd1 _8737__4/HI _8832_/A sky130_fd_sc_hd__conb_1
XFILLER_78_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8811__78 vssd1 vssd1 vccd1 vccd1 _8811__78/HI _8920_/A sky130_fd_sc_hd__conb_1
X_5971_ _5971_/A _6172_/A vssd1 vssd1 vccd1 vccd1 _6194_/B sky130_fd_sc_hd__nand2_1
X_8690_ _8695_/CLK _8690_/D vssd1 vssd1 vccd1 vccd1 _8690_/Q sky130_fd_sc_hd__dfxtp_1
X_4922_ _4937_/A _4990_/B vssd1 vssd1 vccd1 vccd1 _5136_/B sky130_fd_sc_hd__nor2_2
X_7710_ _8515_/C _8124_/A vssd1 vssd1 vccd1 vccd1 _7796_/C sky130_fd_sc_hd__or2_1
X_7641_ _7629_/A _7666_/B _7636_/X _7634_/X vssd1 vssd1 vccd1 vccd1 _7642_/B sky130_fd_sc_hd__a211o_1
XFILLER_33_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4853_ _4879_/A _4906_/A vssd1 vssd1 vccd1 vccd1 _4963_/B sky130_fd_sc_hd__nor2_1
XFILLER_33_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4784_ _4786_/A _4781_/X _4783_/X vssd1 vssd1 vccd1 vccd1 _8620_/D sky130_fd_sc_hd__o21ba_1
X_7572_ _8719_/Q vssd1 vssd1 vccd1 vccd1 _7590_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6523_ _6518_/A _6518_/B _6516_/B vssd1 vssd1 vccd1 vccd1 _6524_/B sky130_fd_sc_hd__a21oi_2
XFILLER_20_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6454_ _6455_/B _6455_/C _6453_/Y vssd1 vssd1 vccd1 vccd1 _8691_/D sky130_fd_sc_hd__a21oi_1
X_5405_ _5404_/B _5426_/B vssd1 vssd1 vccd1 vccd1 _5406_/B sky130_fd_sc_hd__and2b_1
X_6385_ _6437_/B _8683_/Q _6383_/X _6384_/X vssd1 vssd1 vccd1 vccd1 _6385_/X sky130_fd_sc_hd__a31o_1
X_5336_ _6468_/C _5338_/C _5311_/X vssd1 vssd1 vccd1 vccd1 _5336_/Y sky130_fd_sc_hd__o21ai_1
X_8124_ _8124_/A _8321_/B vssd1 vssd1 vccd1 vccd1 _8225_/A sky130_fd_sc_hd__or2_1
X_5267_ _8567_/A vssd1 vssd1 vccd1 vccd1 _5267_/X sky130_fd_sc_hd__clkbuf_2
X_8055_ _8281_/B _8167_/A _8297_/A vssd1 vssd1 vccd1 vccd1 _8087_/B sky130_fd_sc_hd__a21o_1
X_7006_ _7342_/A _7342_/B vssd1 vssd1 vccd1 vccd1 _7015_/A sky130_fd_sc_hd__xnor2_1
XFILLER_87_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5198_ _5195_/X _5196_/X _5197_/X vssd1 vssd1 vccd1 vccd1 _5198_/X sky130_fd_sc_hd__o21a_1
XFILLER_68_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7908_ _7908_/A _8057_/A vssd1 vssd1 vccd1 vccd1 _7910_/A sky130_fd_sc_hd__nor2_1
XFILLER_36_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8888_ _8888_/A _4402_/Y vssd1 vssd1 vccd1 vccd1 io_out[25] sky130_fd_sc_hd__ebufn_8
XFILLER_70_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7839_ _7839_/A _7839_/B vssd1 vssd1 vccd1 vccd1 _8205_/A sky130_fd_sc_hd__nor2_1
Xclkbuf_4_11_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8681_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_50_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6170_ _5976_/A _5976_/B _5974_/Y vssd1 vssd1 vccd1 vccd1 _6177_/A sky130_fd_sc_hd__a21oi_1
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5121_ _5121_/A _5136_/C vssd1 vssd1 vccd1 vccd1 _5230_/D sky130_fd_sc_hd__or2_1
XFILLER_69_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5052_ _4661_/A _5042_/X _5045_/X _4986_/B _5051_/X vssd1 vssd1 vccd1 vccd1 _5052_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_57_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5954_ _6168_/A _5954_/B vssd1 vssd1 vccd1 vccd1 _5955_/B sky130_fd_sc_hd__xnor2_1
X_4905_ _5084_/C _5231_/A vssd1 vssd1 vccd1 vccd1 _4932_/A sky130_fd_sc_hd__or2_1
XFILLER_21_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5885_ _5885_/A vssd1 vssd1 vccd1 vccd1 _6218_/B sky130_fd_sc_hd__clkbuf_2
X_8673_ _8674_/CLK _8673_/D vssd1 vssd1 vccd1 vccd1 _8673_/Q sky130_fd_sc_hd__dfxtp_1
X_4836_ _4839_/A _4848_/A _4848_/B vssd1 vssd1 vccd1 vccd1 _4891_/C sky130_fd_sc_hd__nand3b_4
XFILLER_21_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7624_ _7623_/X _7619_/A _7624_/S vssd1 vssd1 vccd1 vccd1 _7625_/B sky130_fd_sc_hd__mux2_1
X_7555_ _7555_/A vssd1 vssd1 vccd1 vccd1 _7555_/Y sky130_fd_sc_hd__inv_2
X_6506_ _6506_/A vssd1 vssd1 vccd1 vccd1 _8698_/D sky130_fd_sc_hd__clkbuf_1
X_4767_ _4765_/B _4786_/C _4765_/A vssd1 vssd1 vccd1 vccd1 _4768_/C sky130_fd_sc_hd__a21o_1
X_4698_ _5190_/A _4698_/B vssd1 vssd1 vccd1 vccd1 _5064_/A sky130_fd_sc_hd__nand2_2
X_7486_ _7488_/A _7489_/S _7395_/X vssd1 vssd1 vccd1 vccd1 _7486_/Y sky130_fd_sc_hd__a21boi_1
X_6437_ _8686_/Q _6437_/B _6437_/C vssd1 vssd1 vccd1 vccd1 _6441_/B sky130_fd_sc_hd__and3_1
XFILLER_20_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6368_ _8673_/Q _6368_/B vssd1 vssd1 vccd1 vccd1 _6372_/B sky130_fd_sc_hd__nor2_1
X_5319_ _8640_/Q _5322_/C vssd1 vssd1 vccd1 vccd1 _5321_/A sky130_fd_sc_hd__and2_1
XFILLER_88_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8107_ _8098_/A _8098_/B _8106_/X vssd1 vssd1 vccd1 vccd1 _8266_/A sky130_fd_sc_hd__a21o_1
X_6299_ _6299_/A _6299_/B _6299_/C vssd1 vssd1 vccd1 vccd1 _6300_/C sky130_fd_sc_hd__nand3_1
XFILLER_102_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8038_ _8116_/A _8039_/B vssd1 vssd1 vccd1 vccd1 _8040_/A sky130_fd_sc_hd__nor2_1
XFILLER_28_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5670_ _5952_/A vssd1 vssd1 vccd1 vccd1 _6120_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4621_ _4623_/B _4645_/B _4621_/C vssd1 vssd1 vccd1 vccd1 _4622_/A sky130_fd_sc_hd__and3b_1
XFILLER_30_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7340_ _7340_/A _7419_/B vssd1 vssd1 vccd1 vccd1 _7345_/A sky130_fd_sc_hd__xnor2_1
X_4552_ _8630_/Q _4552_/B vssd1 vssd1 vccd1 vccd1 _4553_/A sky130_fd_sc_hd__and2_1
X_7271_ _7272_/A _7272_/B vssd1 vssd1 vccd1 vccd1 _7283_/A sky130_fd_sc_hd__nand2_1
X_4483_ _8621_/Q vssd1 vssd1 vccd1 vccd1 _7906_/B sky130_fd_sc_hd__clkbuf_2
X_6222_ _5901_/A _6004_/A _6221_/X vssd1 vssd1 vccd1 vccd1 _6223_/B sky130_fd_sc_hd__a21o_1
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6153_ _6307_/A _6307_/B vssd1 vssd1 vccd1 vccd1 _6153_/X sky130_fd_sc_hd__or2b_1
X_5104_ _4986_/B _5103_/X _5058_/X vssd1 vssd1 vccd1 vccd1 _5104_/X sky130_fd_sc_hd__a21o_1
XFILLER_85_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6084_ _6084_/A _6141_/A vssd1 vssd1 vccd1 vccd1 _6087_/A sky130_fd_sc_hd__or2b_1
XFILLER_85_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5035_ _5035_/A vssd1 vssd1 vccd1 vccd1 _5208_/A sky130_fd_sc_hd__clkbuf_2
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6986_ _6985_/A _6985_/B _6985_/C vssd1 vssd1 vccd1 vccd1 _6989_/B sky130_fd_sc_hd__a21o_1
XFILLER_80_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8725_ _8735_/CLK _8725_/D vssd1 vssd1 vccd1 vccd1 _8725_/Q sky130_fd_sc_hd__dfxtp_1
X_5937_ _5937_/A _5916_/B vssd1 vssd1 vccd1 vccd1 _5960_/B sky130_fd_sc_hd__or2b_1
X_8656_ _8733_/CLK _8656_/D vssd1 vssd1 vccd1 vccd1 _8656_/Q sky130_fd_sc_hd__dfxtp_1
X_5868_ _5868_/A _5868_/B vssd1 vssd1 vccd1 vccd1 _5869_/B sky130_fd_sc_hd__xnor2_2
X_7607_ _8721_/Q _6423_/X _7606_/X vssd1 vssd1 vccd1 vccd1 _8721_/D sky130_fd_sc_hd__a21bo_1
X_4819_ _4839_/B _4891_/A _4898_/A vssd1 vssd1 vccd1 vccd1 _4863_/A sky130_fd_sc_hd__nor3_1
X_5799_ _5879_/B _5799_/B vssd1 vssd1 vccd1 vccd1 _5800_/B sky130_fd_sc_hd__or2_1
XFILLER_31_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8587_ _8672_/CLK _8587_/D vssd1 vssd1 vccd1 vccd1 _8587_/Q sky130_fd_sc_hd__dfxtp_1
X_7538_ _6508_/A _7547_/S _7536_/Y _7537_/X vssd1 vssd1 vccd1 vccd1 _8713_/D sky130_fd_sc_hd__a31o_1
XFILLER_5_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7469_ _7469_/A _7469_/B vssd1 vssd1 vccd1 vccd1 _7509_/A sky130_fd_sc_hd__xnor2_2
XFILLER_31_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6840_ _6837_/X _7432_/B _7145_/A vssd1 vssd1 vccd1 vccd1 _7072_/A sky130_fd_sc_hd__o21a_1
XFILLER_35_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6771_ _6999_/A _7335_/B vssd1 vssd1 vccd1 vccd1 _7004_/A sky130_fd_sc_hd__xnor2_4
XFILLER_23_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5722_ _5722_/A _5580_/A vssd1 vssd1 vccd1 vccd1 _5722_/X sky130_fd_sc_hd__or2b_1
X_8510_ _8510_/A _8510_/B vssd1 vssd1 vccd1 vccd1 _8510_/Y sky130_fd_sc_hd__nor2_1
X_8441_ _8394_/A _8394_/B _8393_/A vssd1 vssd1 vccd1 vccd1 _8442_/B sky130_fd_sc_hd__a21oi_1
X_5653_ _6028_/A _5910_/B _5820_/A vssd1 vssd1 vccd1 vccd1 _5737_/A sky130_fd_sc_hd__mux2_2
X_8372_ _8372_/A _8372_/B vssd1 vssd1 vccd1 vccd1 _8469_/B sky130_fd_sc_hd__xor2_1
X_5584_ _5584_/A _5584_/B vssd1 vssd1 vccd1 vccd1 _5694_/B sky130_fd_sc_hd__xor2_2
X_4604_ _8586_/Q _8587_/Q _4604_/C vssd1 vssd1 vccd1 vccd1 _4610_/C sky130_fd_sc_hd__and3_1
X_7323_ _6967_/B _6967_/C _6967_/A vssd1 vssd1 vccd1 vccd1 _7340_/A sky130_fd_sc_hd__a21boi_2
X_4535_ _4839_/B vssd1 vssd1 vccd1 vccd1 _4900_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7254_ _7254_/A _7254_/B _7254_/C vssd1 vssd1 vccd1 vccd1 _7256_/A sky130_fd_sc_hd__and3_1
X_4466_ _8609_/Q vssd1 vssd1 vccd1 vccd1 _7677_/B sky130_fd_sc_hd__inv_2
XFILLER_104_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7185_ _7185_/A _7185_/B _7185_/C vssd1 vssd1 vccd1 vccd1 _7188_/A sky130_fd_sc_hd__and3_1
X_4397_ _4400_/A vssd1 vssd1 vccd1 vccd1 _4397_/Y sky130_fd_sc_hd__inv_2
X_6205_ _6118_/A _6020_/Y _6204_/Y vssd1 vssd1 vccd1 vccd1 _6253_/B sky130_fd_sc_hd__a21o_1
X_6136_ _6136_/A _6136_/B vssd1 vssd1 vccd1 vccd1 _6321_/B sky130_fd_sc_hd__nand2_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6067_ _5746_/A _6316_/B _6039_/B _6066_/X vssd1 vssd1 vccd1 vccd1 _6082_/B sky130_fd_sc_hd__a31o_1
X_5018_ _5018_/A vssd1 vssd1 vccd1 vccd1 _5194_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_38_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8772__39 vssd1 vssd1 vccd1 vccd1 _8772__39/HI _8867_/A sky130_fd_sc_hd__conb_1
X_6969_ _7254_/A _7370_/A vssd1 vssd1 vccd1 vccd1 _6975_/A sky130_fd_sc_hd__nor2_1
XFILLER_81_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8708_ _8734_/CLK _8708_/D vssd1 vssd1 vccd1 vccd1 _8708_/Q sky130_fd_sc_hd__dfxtp_1
X_8639_ _8710_/CLK _8639_/D vssd1 vssd1 vccd1 vccd1 _8639_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7941_ _8017_/A _7941_/B vssd1 vssd1 vccd1 vccd1 _8102_/B sky130_fd_sc_hd__or2_2
XFILLER_35_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7872_ _7771_/A _7871_/X _7771_/C _7768_/A vssd1 vssd1 vccd1 vccd1 _7952_/B sky130_fd_sc_hd__a31o_1
XFILLER_63_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6823_ _6927_/A vssd1 vssd1 vccd1 vccd1 _6857_/A sky130_fd_sc_hd__clkinv_2
X_6754_ _7054_/B vssd1 vssd1 vccd1 vccd1 _7196_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_6685_ _6780_/A _6793_/C _6685_/C vssd1 vssd1 vccd1 vccd1 _6697_/A sky130_fd_sc_hd__nand3_1
XFILLER_50_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5705_ _5705_/A _5780_/B _5780_/C vssd1 vssd1 vccd1 vccd1 _5708_/A sky130_fd_sc_hd__and3_2
XFILLER_12_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8424_ _8437_/A _8437_/B vssd1 vssd1 vccd1 vccd1 _8425_/B sky130_fd_sc_hd__xnor2_1
X_5636_ _5811_/A vssd1 vssd1 vccd1 vccd1 _5944_/B sky130_fd_sc_hd__clkbuf_2
X_8355_ _8352_/B _8355_/B vssd1 vssd1 vccd1 vccd1 _8427_/A sky130_fd_sc_hd__and2b_1
X_5567_ _5780_/A _5567_/B vssd1 vssd1 vccd1 vccd1 _6108_/A sky130_fd_sc_hd__nand2_2
X_7306_ _7306_/A _7016_/B vssd1 vssd1 vccd1 vccd1 _7306_/X sky130_fd_sc_hd__or2b_1
X_4518_ _8603_/Q vssd1 vssd1 vccd1 vccd1 _5171_/A sky130_fd_sc_hd__buf_2
X_8286_ _7649_/B _8474_/A _7724_/Y vssd1 vssd1 vccd1 vccd1 _8365_/C sky130_fd_sc_hd__o21a_1
X_5498_ _5498_/A _5575_/A vssd1 vssd1 vccd1 vccd1 _5539_/C sky130_fd_sc_hd__xnor2_1
X_4449_ _4449_/A vssd1 vssd1 vccd1 vccd1 _4449_/Y sky130_fd_sc_hd__inv_2
X_7237_ _7454_/A _7172_/C _7236_/X vssd1 vssd1 vccd1 vccd1 _7238_/B sky130_fd_sc_hd__a21oi_2
X_8817__84 vssd1 vssd1 vccd1 vccd1 _8817__84/HI _8926_/A sky130_fd_sc_hd__conb_1
X_7168_ _7212_/A _7212_/B vssd1 vssd1 vccd1 vccd1 _7187_/A sky130_fd_sc_hd__nor2_1
X_7099_ _7099_/A _7099_/B _7099_/C vssd1 vssd1 vccd1 vccd1 _7124_/D sky130_fd_sc_hd__nand3_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6119_ _6119_/A _6119_/B vssd1 vssd1 vccd1 vccd1 _6120_/B sky130_fd_sc_hd__nand2_1
XFILLER_100_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6470_ _8649_/Q _8648_/Q _8653_/Q _8652_/Q vssd1 vssd1 vccd1 vccd1 _6471_/D sky130_fd_sc_hd__and4_1
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5421_ _5420_/X _5415_/B _5413_/B vssd1 vssd1 vccd1 vccd1 _5423_/C sky130_fd_sc_hd__a21oi_1
X_5352_ _8650_/Q _5350_/A _5311_/X vssd1 vssd1 vccd1 vccd1 _5353_/B sky130_fd_sc_hd__o21ai_1
X_8140_ _8139_/B _8321_/B _8450_/B vssd1 vssd1 vccd1 vccd1 _8402_/A sky130_fd_sc_hd__a21o_2
XFILLER_99_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8071_ _8071_/A _8368_/A vssd1 vssd1 vccd1 vccd1 _8072_/D sky130_fd_sc_hd__or2b_1
X_7022_ _7039_/A vssd1 vssd1 vccd1 vccd1 _7403_/A sky130_fd_sc_hd__clkbuf_2
X_5283_ _8632_/Q _5285_/B vssd1 vssd1 vccd1 vccd1 _5283_/X sky130_fd_sc_hd__or2_1
XINSDIODE2_9 _4928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7924_ _7819_/A _7819_/B _7923_/Y vssd1 vssd1 vccd1 vccd1 _7926_/B sky130_fd_sc_hd__a21oi_1
XFILLER_43_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7855_ _7792_/A _7792_/B _7854_/X vssd1 vssd1 vccd1 vccd1 _7946_/A sky130_fd_sc_hd__a21o_1
X_6806_ _6806_/A _6806_/B vssd1 vssd1 vccd1 vccd1 _6816_/A sky130_fd_sc_hd__xnor2_1
XFILLER_11_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4998_ _5244_/B _4998_/B _5091_/C vssd1 vssd1 vccd1 vccd1 _5236_/C sky130_fd_sc_hd__or3_1
XFILLER_51_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7786_ _7950_/A vssd1 vssd1 vccd1 vccd1 _7960_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_23_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6737_ _6715_/A _7130_/A _7133_/A _7088_/B vssd1 vssd1 vccd1 vccd1 _7076_/B sky130_fd_sc_hd__a22o_1
XFILLER_23_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6668_ _7075_/A _7074_/B _7074_/C _6972_/C _7350_/B vssd1 vssd1 vccd1 vccd1 _6669_/A
+ sky130_fd_sc_hd__o32ai_2
X_6599_ _8609_/Q _8713_/Q vssd1 vssd1 vccd1 vccd1 _6826_/A sky130_fd_sc_hd__or2b_2
X_8407_ _8407_/A _8407_/B vssd1 vssd1 vccd1 vccd1 _8443_/A sky130_fd_sc_hd__xnor2_2
X_5619_ _5619_/A _5619_/B vssd1 vssd1 vccd1 vccd1 _5630_/A sky130_fd_sc_hd__nand2_2
X_8338_ _8338_/A _8338_/B vssd1 vssd1 vccd1 vccd1 _8415_/C sky130_fd_sc_hd__xnor2_1
XFILLER_2_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8269_ _8269_/A _8269_/B vssd1 vssd1 vccd1 vccd1 _8501_/B sky130_fd_sc_hd__nor2_1
XFILLER_59_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5970_ _5970_/A _5970_/B vssd1 vssd1 vccd1 vccd1 _5974_/B sky130_fd_sc_hd__nand2_1
XFILLER_25_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4921_ _5007_/A _4963_/B _5173_/B vssd1 vssd1 vccd1 vccd1 _5210_/B sky130_fd_sc_hd__or3b_2
X_4852_ _4852_/A _5087_/A vssd1 vssd1 vccd1 vccd1 _4906_/A sky130_fd_sc_hd__nor2_2
X_7640_ _7834_/A vssd1 vssd1 vccd1 vccd1 _8066_/A sky130_fd_sc_hd__clkinv_2
X_4783_ _4786_/A _4790_/A _4779_/B _4785_/A vssd1 vssd1 vccd1 vccd1 _4783_/X sky130_fd_sc_hd__a31o_1
X_7571_ _7596_/B _8717_/Q vssd1 vssd1 vccd1 vccd1 _7597_/A sky130_fd_sc_hd__and2b_1
X_6522_ _6520_/Y _6522_/B vssd1 vssd1 vccd1 vccd1 _6524_/A sky130_fd_sc_hd__and2b_1
X_6453_ _6455_/B _6455_/C _6401_/B vssd1 vssd1 vccd1 vccd1 _6453_/Y sky130_fd_sc_hd__o21ai_1
X_5404_ _8656_/Q _5404_/B vssd1 vssd1 vccd1 vccd1 _5406_/A sky130_fd_sc_hd__and2b_1
X_6384_ _8685_/Q _8684_/Q _8686_/Q vssd1 vssd1 vccd1 vccd1 _6384_/X sky130_fd_sc_hd__a21o_1
X_8123_ _8399_/B _8229_/A _8123_/S vssd1 vssd1 vccd1 vccd1 _8323_/A sky130_fd_sc_hd__mux2_1
X_5335_ _8645_/Q vssd1 vssd1 vccd1 vccd1 _6468_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_87_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5266_ _8625_/Q _5276_/B vssd1 vssd1 vccd1 vccd1 _5266_/X sky130_fd_sc_hd__or2_1
X_8054_ _8054_/A _8365_/B vssd1 vssd1 vccd1 vccd1 _8297_/A sky130_fd_sc_hd__nand2_1
XFILLER_102_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7005_ _6911_/A _6911_/B _7004_/X vssd1 vssd1 vccd1 vccd1 _7342_/B sky130_fd_sc_hd__a21oi_1
X_5197_ _4923_/X _5238_/C _5170_/B _5059_/X _5069_/X vssd1 vssd1 vccd1 vccd1 _5197_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_95_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7907_ _7802_/B _7804_/B _7906_/X vssd1 vssd1 vccd1 vccd1 _8057_/A sky130_fd_sc_hd__a21o_1
X_8887_ _8887_/A _4400_/Y vssd1 vssd1 vccd1 vccd1 io_out[24] sky130_fd_sc_hd__ebufn_8
XFILLER_24_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7838_ _8208_/A _8139_/A vssd1 vssd1 vccd1 vccd1 _7839_/B sky130_fd_sc_hd__nor2_1
X_7769_ _7769_/A _7769_/B vssd1 vssd1 vccd1 vccd1 _7769_/X sky130_fd_sc_hd__or2_1
XFILLER_11_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5120_ _5120_/A _5120_/B _5227_/C _5120_/D vssd1 vssd1 vccd1 vccd1 _5120_/X sky130_fd_sc_hd__or4_1
XFILLER_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5051_ _5215_/A _5078_/C _5200_/C _5050_/X _5009_/B vssd1 vssd1 vccd1 vccd1 _5051_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_57_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5953_ _5953_/A _5953_/B _6171_/B vssd1 vssd1 vccd1 vccd1 _5954_/B sky130_fd_sc_hd__and3_1
X_4904_ _4904_/A _4904_/B vssd1 vssd1 vccd1 vccd1 _5231_/A sky130_fd_sc_hd__nor2_2
X_8672_ _8672_/CLK _8672_/D vssd1 vssd1 vccd1 vccd1 _8672_/Q sky130_fd_sc_hd__dfxtp_1
X_5884_ _6204_/A _5884_/B vssd1 vssd1 vccd1 vccd1 _5885_/A sky130_fd_sc_hd__nor2_1
XFILLER_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4835_ _4948_/B _4837_/B vssd1 vssd1 vccd1 vccd1 _4955_/A sky130_fd_sc_hd__nor2_1
X_7623_ _8722_/Q _7623_/B vssd1 vssd1 vccd1 vccd1 _7623_/X sky130_fd_sc_hd__or2_1
X_4766_ _4774_/C vssd1 vssd1 vccd1 vccd1 _4779_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_21_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7554_ _8735_/Q vssd1 vssd1 vccd1 vccd1 _7876_/A sky130_fd_sc_hd__clkbuf_2
X_6505_ _5362_/A _6507_/A _6565_/A vssd1 vssd1 vccd1 vccd1 _6506_/A sky130_fd_sc_hd__mux2_1
X_4697_ _5065_/A vssd1 vssd1 vccd1 vccd1 _4697_/X sky130_fd_sc_hd__clkbuf_2
X_7485_ _7475_/X _7476_/Y _7480_/X _7482_/Y _7484_/Y vssd1 vssd1 vccd1 vccd1 _7491_/C
+ sky130_fd_sc_hd__o2111a_1
XFILLER_20_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6436_ _6437_/B _6437_/C _6435_/Y vssd1 vssd1 vccd1 vccd1 _8685_/D sky130_fd_sc_hd__a21oi_1
XFILLER_20_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6367_ _8673_/Q _6368_/B vssd1 vssd1 vccd1 vccd1 _6369_/A sky130_fd_sc_hd__and2_1
X_5318_ _5318_/A vssd1 vssd1 vccd1 vccd1 _8639_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8106_ _8097_/B _8106_/B vssd1 vssd1 vccd1 vccd1 _8106_/X sky130_fd_sc_hd__and2b_1
XFILLER_102_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6298_ _6298_/A _6298_/B vssd1 vssd1 vccd1 vccd1 _6332_/A sky130_fd_sc_hd__and2_1
XFILLER_102_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5249_ _5079_/A _5212_/B _5242_/X _5248_/X _5080_/Y vssd1 vssd1 vccd1 vccd1 _5249_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8037_ _8217_/A _7960_/B _7965_/B _7963_/X vssd1 vssd1 vccd1 vccd1 _8039_/B sky130_fd_sc_hd__a31oi_1
XFILLER_75_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8778__45 vssd1 vssd1 vccd1 vccd1 _8778__45/HI _8873_/A sky130_fd_sc_hd__conb_1
XFILLER_19_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4620_ _8590_/Q _8591_/Q _4614_/B _8592_/Q vssd1 vssd1 vccd1 vccd1 _4621_/C sky130_fd_sc_hd__a31o_1
X_4551_ _4551_/A vssd1 vssd1 vccd1 vccd1 _8879_/A sky130_fd_sc_hd__clkbuf_1
X_4482_ _4482_/A vssd1 vssd1 vccd1 vccd1 _8874_/A sky130_fd_sc_hd__clkbuf_1
X_7270_ _7270_/A _7270_/B vssd1 vssd1 vccd1 vccd1 _7283_/B sky130_fd_sc_hd__xor2_2
X_6221_ _6221_/A _6221_/B _6221_/C vssd1 vssd1 vccd1 vccd1 _6221_/X sky130_fd_sc_hd__and3_1
XFILLER_103_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6152_ _6152_/A _6152_/B vssd1 vssd1 vccd1 vccd1 _6307_/B sky130_fd_sc_hd__xor2_1
X_5103_ _5103_/A _5103_/B vssd1 vssd1 vccd1 vccd1 _5103_/X sky130_fd_sc_hd__or2_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6083_ _6084_/A _6083_/B _6083_/C vssd1 vssd1 vccd1 vccd1 _6141_/A sky130_fd_sc_hd__or3_1
XFILLER_85_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5034_ _6603_/B _5034_/B vssd1 vssd1 vccd1 vccd1 _5256_/A sky130_fd_sc_hd__xnor2_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6985_ _6985_/A _6985_/B _6985_/C vssd1 vssd1 vccd1 vccd1 _6989_/A sky130_fd_sc_hd__nand3_1
XFILLER_53_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5936_ _5936_/A _5936_/B vssd1 vssd1 vccd1 vccd1 _5960_/A sky130_fd_sc_hd__nand2_1
XFILLER_15_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8724_ _8735_/CLK _8724_/D vssd1 vssd1 vccd1 vccd1 _8724_/Q sky130_fd_sc_hd__dfxtp_1
X_8655_ _8671_/CLK _8655_/D vssd1 vssd1 vccd1 vccd1 _8655_/Q sky130_fd_sc_hd__dfxtp_1
X_5867_ _5979_/A _5867_/B vssd1 vssd1 vccd1 vccd1 _5868_/B sky130_fd_sc_hd__or2_1
XFILLER_21_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7606_ _7603_/X _7604_/X _7605_/Y _8578_/A vssd1 vssd1 vccd1 vccd1 _7606_/X sky130_fd_sc_hd__a211o_1
X_4818_ _4898_/A _4818_/B vssd1 vssd1 vccd1 vccd1 _5066_/A sky130_fd_sc_hd__nor2_1
XFILLER_21_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5798_ _5798_/A _5798_/B vssd1 vssd1 vccd1 vccd1 _5799_/B sky130_fd_sc_hd__nor2_1
X_8586_ _8672_/CLK _8586_/D vssd1 vssd1 vccd1 vccd1 _8586_/Q sky130_fd_sc_hd__dfxtp_1
X_7537_ _7546_/A _7537_/B _7537_/C vssd1 vssd1 vccd1 vccd1 _7537_/X sky130_fd_sc_hd__and3_1
X_4749_ _4749_/A _4900_/A _4957_/A vssd1 vssd1 vccd1 vccd1 _4758_/B sky130_fd_sc_hd__and3_1
X_7468_ _7468_/A _7468_/B vssd1 vssd1 vccd1 vccd1 _7491_/A sky130_fd_sc_hd__xnor2_2
X_6419_ _8678_/Q _6394_/D _6413_/B _8680_/Q vssd1 vssd1 vccd1 vccd1 _6420_/B sky130_fd_sc_hd__a31o_1
X_7399_ _7399_/A _7392_/A vssd1 vssd1 vccd1 vccd1 _7399_/X sky130_fd_sc_hd__or2b_1
XFILLER_103_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6770_ _7409_/A _6713_/B vssd1 vssd1 vccd1 vccd1 _6868_/A sky130_fd_sc_hd__or2b_1
XFILLER_50_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5721_ _5721_/A _5721_/B vssd1 vssd1 vccd1 vccd1 _5726_/A sky130_fd_sc_hd__xor2_2
X_8440_ _8382_/A _8382_/B _8439_/X vssd1 vssd1 vccd1 vccd1 _8467_/A sky130_fd_sc_hd__a21oi_1
X_5652_ _5652_/A _5811_/A vssd1 vssd1 vccd1 vccd1 _5820_/A sky130_fd_sc_hd__nand2_1
XFILLER_30_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8371_ _8371_/A _8471_/B vssd1 vssd1 vccd1 vccd1 _8372_/B sky130_fd_sc_hd__xnor2_1
X_5583_ _5583_/A _5696_/B vssd1 vssd1 vccd1 vccd1 _5584_/B sky130_fd_sc_hd__xnor2_2
XFILLER_30_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4603_ _4603_/A _4603_/B vssd1 vssd1 vccd1 vccd1 _8586_/D sky130_fd_sc_hd__nor2_1
X_7322_ _7322_/A _7322_/B vssd1 vssd1 vccd1 vccd1 _7388_/A sky130_fd_sc_hd__xnor2_1
X_4534_ _4845_/C vssd1 vssd1 vccd1 vccd1 _4839_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4465_ _8610_/Q vssd1 vssd1 vccd1 vccd1 _6605_/B sky130_fd_sc_hd__clkbuf_2
X_7253_ _7335_/A _7261_/B vssd1 vssd1 vccd1 vccd1 _7274_/A sky130_fd_sc_hd__xnor2_2
X_7184_ _7143_/B _7143_/C _7143_/A vssd1 vssd1 vccd1 vccd1 _7185_/C sky130_fd_sc_hd__a21o_1
X_4396_ _4400_/A vssd1 vssd1 vccd1 vccd1 _4396_/Y sky130_fd_sc_hd__inv_2
X_6204_ _6204_/A _6204_/B vssd1 vssd1 vccd1 vccd1 _6204_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_58_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6135_ _6126_/A _6126_/C _6126_/B vssd1 vssd1 vccd1 vccd1 _6136_/B sky130_fd_sc_hd__o21ai_1
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6066_ _6038_/A _6066_/B vssd1 vssd1 vccd1 vccd1 _6066_/X sky130_fd_sc_hd__and2b_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5017_ _5215_/A _5154_/A _5017_/C _5153_/B vssd1 vssd1 vccd1 vccd1 _5017_/X sky130_fd_sc_hd__or4_1
XFILLER_53_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6968_ _6967_/A _6967_/B _6967_/C vssd1 vssd1 vccd1 vccd1 _7347_/B sky130_fd_sc_hd__a21oi_1
X_8707_ _8734_/CLK _8707_/D vssd1 vssd1 vccd1 vccd1 _8707_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6899_ _6952_/A _6952_/B vssd1 vssd1 vccd1 vccd1 _6901_/C sky130_fd_sc_hd__xnor2_2
X_5919_ _5919_/A _5919_/B vssd1 vssd1 vccd1 vccd1 _5920_/B sky130_fd_sc_hd__nand2_1
X_8638_ _8710_/CLK _8638_/D vssd1 vssd1 vccd1 vccd1 _8638_/Q sky130_fd_sc_hd__dfxtp_1
X_8569_ _8569_/A _8577_/S vssd1 vssd1 vccd1 vccd1 _8573_/A sky130_fd_sc_hd__or2b_1
XFILLER_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8748__15 vssd1 vssd1 vccd1 vccd1 _8748__15/HI _8843_/A sky130_fd_sc_hd__conb_1
XFILLER_76_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7940_ _7940_/A _7940_/B _7940_/C vssd1 vssd1 vccd1 vccd1 _7941_/B sky130_fd_sc_hd__and3_1
X_7871_ _7871_/A _8735_/Q vssd1 vssd1 vccd1 vccd1 _7871_/X sky130_fd_sc_hd__or2b_1
X_6822_ _6841_/A vssd1 vssd1 vccd1 vccd1 _7409_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_90_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6753_ _7063_/B vssd1 vssd1 vccd1 vccd1 _6841_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_50_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6684_ _6669_/A _6672_/A _6715_/A vssd1 vssd1 vccd1 vccd1 _6685_/C sky130_fd_sc_hd__a21o_1
X_5704_ _5781_/A vssd1 vssd1 vccd1 vccd1 _5987_/A sky130_fd_sc_hd__buf_2
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8423_ _8423_/A _8487_/B vssd1 vssd1 vccd1 vccd1 _8437_/B sky130_fd_sc_hd__xnor2_1
X_5635_ _5609_/B _5614_/B _5634_/X vssd1 vssd1 vccd1 vccd1 _5811_/A sky130_fd_sc_hd__a21oi_1
XFILLER_31_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8354_ _8431_/A _8431_/B vssd1 vssd1 vccd1 vccd1 _8429_/A sky130_fd_sc_hd__nand2_1
X_5566_ _5566_/A vssd1 vssd1 vccd1 vccd1 _6204_/A sky130_fd_sc_hd__clkbuf_2
X_7305_ _7403_/A _7303_/Y _7304_/Y vssd1 vssd1 vccd1 vccd1 _7322_/A sky130_fd_sc_hd__a21o_1
X_4517_ _4986_/A vssd1 vssd1 vccd1 vccd1 _5190_/A sky130_fd_sc_hd__clkbuf_2
X_8285_ _8284_/A _8367_/A _8291_/B _8291_/A vssd1 vssd1 vccd1 vccd1 _8289_/A sky130_fd_sc_hd__o22ai_2
X_5497_ _5502_/A _5780_/B _5780_/C vssd1 vssd1 vccd1 vccd1 _5575_/A sky130_fd_sc_hd__and3_2
XFILLER_104_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4448_ _4449_/A vssd1 vssd1 vccd1 vccd1 _4448_/Y sky130_fd_sc_hd__inv_2
X_7236_ _7128_/A _7213_/B _7254_/C _6711_/A vssd1 vssd1 vccd1 vccd1 _7236_/X sky130_fd_sc_hd__o22a_1
XFILLER_104_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4379_ _4382_/A vssd1 vssd1 vccd1 vccd1 _4379_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7167_ _7167_/A _7167_/B vssd1 vssd1 vccd1 vccd1 _7212_/B sky130_fd_sc_hd__or2_1
XFILLER_100_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7098_ _7151_/A _7151_/B _7112_/B _7097_/B _7097_/A vssd1 vssd1 vccd1 vccd1 _7162_/A
+ sky130_fd_sc_hd__a32o_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6118_ _6118_/A _6134_/A vssd1 vssd1 vccd1 vccd1 _6126_/A sky130_fd_sc_hd__nor2_1
XFILLER_85_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6049_ _6049_/A _6049_/B vssd1 vssd1 vccd1 vccd1 _6049_/Y sky130_fd_sc_hd__nor2_1
XFILLER_39_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5420_ _5426_/B _5411_/B vssd1 vssd1 vccd1 vccd1 _5420_/X sky130_fd_sc_hd__or2b_1
X_5351_ _8649_/Q _8650_/Q _5351_/C vssd1 vssd1 vccd1 vccd1 _5354_/B sky130_fd_sc_hd__and3_1
X_5282_ _8706_/Q _5271_/X _5281_/X _5279_/X vssd1 vssd1 vccd1 vccd1 _8631_/D sky130_fd_sc_hd__o211a_1
X_8070_ _8304_/A vssd1 vssd1 vccd1 vccd1 _8368_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7021_ _7018_/Y _7019_/X _6902_/A _6950_/X vssd1 vssd1 vccd1 vccd1 _7042_/B sky130_fd_sc_hd__o211a_1
XFILLER_101_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7923_ _7923_/A _7923_/B vssd1 vssd1 vccd1 vccd1 _7923_/Y sky130_fd_sc_hd__nor2_1
XFILLER_82_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7854_ _8203_/A _8515_/D _7854_/C vssd1 vssd1 vccd1 vccd1 _7854_/X sky130_fd_sc_hd__and3_1
X_6805_ _6803_/X _7103_/A _6804_/X vssd1 vssd1 vccd1 vccd1 _6806_/B sky130_fd_sc_hd__o21ba_1
XFILLER_51_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7785_ _7785_/A vssd1 vssd1 vccd1 vccd1 _7950_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4997_ _5016_/A _5192_/A vssd1 vssd1 vccd1 vccd1 _5155_/C sky130_fd_sc_hd__or2_1
X_6736_ _6972_/C _7080_/A vssd1 vssd1 vccd1 vccd1 _7088_/B sky130_fd_sc_hd__xnor2_2
XFILLER_51_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6667_ _6734_/B vssd1 vssd1 vccd1 vccd1 _7350_/B sky130_fd_sc_hd__clkbuf_2
X_6598_ _6598_/A _8714_/Q vssd1 vssd1 vccd1 vccd1 _6825_/A sky130_fd_sc_hd__or2b_1
X_5618_ _5642_/A _5638_/B vssd1 vssd1 vccd1 vccd1 _5952_/A sky130_fd_sc_hd__xnor2_4
X_8406_ _8325_/A _8325_/B _8324_/A vssd1 vssd1 vccd1 vccd1 _8407_/B sky130_fd_sc_hd__a21oi_2
XFILLER_3_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5549_ _5584_/A _5549_/B vssd1 vssd1 vccd1 vccd1 _5549_/Y sky130_fd_sc_hd__nor2_1
X_8337_ _8397_/B _8337_/B vssd1 vssd1 vccd1 vccd1 _8343_/A sky130_fd_sc_hd__xnor2_1
X_8268_ _8509_/B _8509_/C _8264_/Y _8509_/A vssd1 vssd1 vccd1 vccd1 _8496_/B sky130_fd_sc_hd__a211o_1
XFILLER_78_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7219_ _7220_/A _7220_/B vssd1 vssd1 vccd1 vccd1 _7219_/Y sky130_fd_sc_hd__nor2_1
X_8199_ _8199_/A _8199_/B vssd1 vssd1 vccd1 vccd1 _8200_/B sky130_fd_sc_hd__xnor2_1
XFILLER_58_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_3_6_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_6_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_65_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4920_ _4937_/A _4920_/B vssd1 vssd1 vccd1 vccd1 _5173_/B sky130_fd_sc_hd__or2_2
XFILLER_64_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4851_ _5047_/A vssd1 vssd1 vccd1 vccd1 _4852_/A sky130_fd_sc_hd__inv_2
XFILLER_33_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4782_ _6503_/A vssd1 vssd1 vccd1 vccd1 _4785_/A sky130_fd_sc_hd__buf_2
XFILLER_20_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7570_ _8720_/Q vssd1 vssd1 vccd1 vccd1 _7596_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6521_ _6521_/A _6526_/B vssd1 vssd1 vccd1 vccd1 _6522_/B sky130_fd_sc_hd__nand2_1
X_6452_ _6455_/C _6452_/B vssd1 vssd1 vccd1 vccd1 _8690_/D sky130_fd_sc_hd__nor2_1
XFILLER_9_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5403_ _5400_/A _5397_/X _5398_/X _5402_/Y vssd1 vssd1 vccd1 vccd1 _8658_/D sky130_fd_sc_hd__a22o_1
X_6383_ _6426_/A _8680_/Q _6382_/X _8682_/Q vssd1 vssd1 vccd1 vccd1 _6383_/X sky130_fd_sc_hd__a211o_1
X_8122_ _8204_/A _8122_/B _8122_/C vssd1 vssd1 vccd1 vccd1 _8229_/A sky130_fd_sc_hd__and3b_1
X_5334_ _5338_/C _5334_/B vssd1 vssd1 vccd1 vccd1 _8644_/D sky130_fd_sc_hd__nor2_1
X_5265_ _5265_/A vssd1 vssd1 vccd1 vccd1 _5276_/B sky130_fd_sc_hd__clkbuf_2
X_8053_ _8146_/B vssd1 vssd1 vccd1 vccd1 _8365_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_7004_ _7004_/A _7327_/A vssd1 vssd1 vccd1 vccd1 _7004_/X sky130_fd_sc_hd__and2_1
XFILLER_87_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5196_ _5226_/B _5196_/B _5207_/A _5218_/A vssd1 vssd1 vccd1 vccd1 _5196_/X sky130_fd_sc_hd__or4_1
XFILLER_18_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8802__69 vssd1 vssd1 vccd1 vccd1 _8802__69/HI _8911_/A sky130_fd_sc_hd__conb_1
XFILLER_55_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8886_ _8886_/A _4399_/Y vssd1 vssd1 vccd1 vccd1 io_out[23] sky130_fd_sc_hd__ebufn_8
X_7906_ _7577_/X _7906_/B vssd1 vssd1 vccd1 vccd1 _7906_/X sky130_fd_sc_hd__and2b_1
XFILLER_36_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7837_ _7859_/B vssd1 vssd1 vccd1 vccd1 _8208_/A sky130_fd_sc_hd__clkbuf_2
X_7768_ _7768_/A _7768_/B vssd1 vssd1 vccd1 vccd1 _7771_/B sky130_fd_sc_hd__nor2_1
X_6719_ _6716_/X _6780_/A _6780_/B vssd1 vssd1 vccd1 vccd1 _6725_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7699_ _7711_/A _7711_/B vssd1 vssd1 vccd1 vccd1 _7758_/A sky130_fd_sc_hd__xor2_1
XFILLER_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5050_ _5207_/B _5229_/B _5050_/C vssd1 vssd1 vccd1 vccd1 _5050_/X sky130_fd_sc_hd__or3_1
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5952_ _5952_/A _5952_/B _5952_/C _5947_/X vssd1 vssd1 vccd1 vccd1 _6171_/B sky130_fd_sc_hd__or4b_1
XFILLER_80_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4903_ _4937_/B _4903_/B vssd1 vssd1 vccd1 vccd1 _5084_/C sky130_fd_sc_hd__nor2_2
XFILLER_52_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8671_ _8671_/CLK _8671_/D vssd1 vssd1 vccd1 vccd1 _8671_/Q sky130_fd_sc_hd__dfxtp_1
X_5883_ _5881_/X _5800_/B _5882_/X vssd1 vssd1 vccd1 vccd1 _5904_/A sky130_fd_sc_hd__o21bai_2
XFILLER_33_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4834_ _4845_/B _4845_/C _4834_/C _4845_/A vssd1 vssd1 vccd1 vccd1 _4948_/B sky130_fd_sc_hd__or4b_4
X_7622_ _7618_/A _7584_/X _7621_/Y _7544_/X vssd1 vssd1 vccd1 vccd1 _8723_/D sky130_fd_sc_hd__a211o_1
X_4765_ _4765_/A _4765_/B _4786_/C vssd1 vssd1 vccd1 vccd1 _4774_/C sky130_fd_sc_hd__and3_1
X_7553_ _8733_/Q vssd1 vssd1 vccd1 vccd1 _8576_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6504_ _8698_/Q vssd1 vssd1 vccd1 vccd1 _6565_/A sky130_fd_sc_hd__inv_2
X_4696_ _5079_/A vssd1 vssd1 vccd1 vccd1 _5065_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7484_ _7484_/A _7484_/B vssd1 vssd1 vccd1 vccd1 _7484_/Y sky130_fd_sc_hd__xnor2_1
X_6435_ _6437_/B _6437_/C _6401_/B vssd1 vssd1 vccd1 vccd1 _6435_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6366_ _6366_/A _6373_/S vssd1 vssd1 vccd1 vccd1 _6370_/A sky130_fd_sc_hd__nand2_1
XFILLER_102_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5317_ _5322_/C _5317_/B _5362_/A vssd1 vssd1 vccd1 vccd1 _5318_/A sky130_fd_sc_hd__and3b_1
X_8105_ _8503_/A _8506_/B _8503_/B vssd1 vssd1 vccd1 vccd1 _8509_/C sky130_fd_sc_hd__a21bo_1
XFILLER_88_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6297_ _6297_/A _6322_/A vssd1 vssd1 vccd1 vccd1 _6298_/B sky130_fd_sc_hd__or2_1
X_8036_ _7972_/A _8321_/B _7973_/B _8325_/A vssd1 vssd1 vccd1 vccd1 _8041_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_88_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5248_ _5248_/A _5248_/B _5248_/C vssd1 vssd1 vccd1 vccd1 _5248_/X sky130_fd_sc_hd__or3_1
XFILLER_29_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5179_ _5230_/A _5179_/B vssd1 vssd1 vccd1 vccd1 _5179_/X sky130_fd_sc_hd__or2_1
XFILLER_75_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8938_ _8938_/A _4460_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[37] sky130_fd_sc_hd__ebufn_8
XFILLER_45_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8869_ _8869_/A _4379_/Y vssd1 vssd1 vccd1 vccd1 io_out[6] sky130_fd_sc_hd__ebufn_8
XFILLER_51_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4550_ _8625_/Q _4552_/B vssd1 vssd1 vccd1 vccd1 _4551_/A sky130_fd_sc_hd__and2_1
X_4481_ _4541_/A _4718_/A vssd1 vssd1 vccd1 vccd1 _4482_/A sky130_fd_sc_hd__or2_1
XFILLER_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6220_ _6220_/A _6220_/B vssd1 vssd1 vccd1 vccd1 _6223_/A sky130_fd_sc_hd__xor2_2
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6151_ _6151_/A _6154_/D vssd1 vssd1 vccd1 vccd1 _6307_/A sky130_fd_sc_hd__and2_1
X_5102_ _5139_/D _5102_/B vssd1 vssd1 vccd1 vccd1 _5103_/B sky130_fd_sc_hd__or2_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6082_ _6082_/A _6082_/B vssd1 vssd1 vccd1 vccd1 _6083_/C sky130_fd_sc_hd__xor2_1
XFILLER_97_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5033_ _6603_/B _6746_/B _5149_/S _5032_/X vssd1 vssd1 vccd1 vccd1 _5033_/X sky130_fd_sc_hd__or4b_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6984_ _6984_/A _6984_/B vssd1 vssd1 vccd1 vccd1 _6985_/C sky130_fd_sc_hd__xor2_1
XFILLER_53_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5935_ _5868_/A _5868_/B _5869_/B _5869_/A vssd1 vssd1 vccd1 vccd1 _5963_/A sky130_fd_sc_hd__o22a_1
XFILLER_15_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8723_ _8732_/CLK _8723_/D vssd1 vssd1 vccd1 vccd1 _8723_/Q sky130_fd_sc_hd__dfxtp_1
X_8654_ _8677_/CLK _8654_/D vssd1 vssd1 vccd1 vccd1 _8654_/Q sky130_fd_sc_hd__dfxtp_1
X_5866_ _6196_/A _5866_/B vssd1 vssd1 vccd1 vccd1 _5867_/B sky130_fd_sc_hd__nor2_1
X_4817_ _5111_/B vssd1 vssd1 vccd1 vccd1 _5188_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_21_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7605_ _7603_/X _7604_/X _7499_/A vssd1 vssd1 vccd1 vccd1 _7605_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_21_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5797_ _5798_/A _5798_/B vssd1 vssd1 vccd1 vccd1 _5879_/B sky130_fd_sc_hd__and2_1
XFILLER_31_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8585_ _8672_/CLK _8585_/D vssd1 vssd1 vccd1 vccd1 _8585_/Q sky130_fd_sc_hd__dfxtp_1
X_7536_ _7535_/A _7535_/C _7535_/B vssd1 vssd1 vccd1 vccd1 _7536_/Y sky130_fd_sc_hd__o21ai_1
X_4748_ _5296_/A vssd1 vssd1 vccd1 vccd1 _7550_/A sky130_fd_sc_hd__clkbuf_2
X_7467_ _7467_/A _7467_/B vssd1 vssd1 vccd1 vccd1 _7468_/B sky130_fd_sc_hd__xnor2_2
X_4679_ _4702_/A _4702_/B vssd1 vssd1 vccd1 vccd1 _4689_/B sky130_fd_sc_hd__nand2_1
X_6418_ _8679_/Q _8680_/Q _6418_/C vssd1 vssd1 vccd1 vccd1 _6426_/C sky130_fd_sc_hd__and3_1
X_7398_ _7488_/A _7489_/S _7394_/X _7396_/X _7397_/X vssd1 vssd1 vccd1 vccd1 _7468_/A
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6349_ _6350_/A _6350_/B vssd1 vssd1 vccd1 vccd1 _6355_/B sky130_fd_sc_hd__or2_1
XFILLER_88_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8019_ _8019_/A _8017_/B vssd1 vssd1 vccd1 vccd1 _8265_/A sky130_fd_sc_hd__or2b_1
XFILLER_56_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5720_ _5720_/A _5720_/B vssd1 vssd1 vccd1 vccd1 _5721_/B sky130_fd_sc_hd__xnor2_1
XFILLER_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5651_ _5746_/A _5859_/B vssd1 vssd1 vccd1 vccd1 _5833_/A sky130_fd_sc_hd__nand2_2
XFILLER_30_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8370_ _8370_/A _8370_/B vssd1 vssd1 vccd1 vccd1 _8471_/B sky130_fd_sc_hd__xnor2_1
X_5582_ _5582_/A _5582_/B vssd1 vssd1 vccd1 vccd1 _5696_/B sky130_fd_sc_hd__xnor2_1
X_4602_ _8586_/Q _4604_/C _4595_/X vssd1 vssd1 vccd1 vccd1 _4603_/B sky130_fd_sc_hd__o21ai_1
X_7321_ _7406_/B _7321_/B vssd1 vssd1 vccd1 vccd1 _7322_/B sky130_fd_sc_hd__xnor2_1
X_4533_ _8613_/Q vssd1 vssd1 vccd1 vccd1 _4845_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_7252_ _7252_/A _7252_/B vssd1 vssd1 vccd1 vccd1 _7264_/A sky130_fd_sc_hd__xor2_2
XFILLER_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6203_ _6000_/A _6000_/B _6202_/X vssd1 vssd1 vccd1 vccd1 _6239_/A sky130_fd_sc_hd__a21o_1
X_4464_ _4464_/A vssd1 vssd1 vccd1 vccd1 _4464_/Y sky130_fd_sc_hd__inv_2
X_7183_ _7208_/A _7208_/B vssd1 vssd1 vccd1 vccd1 _7185_/B sky130_fd_sc_hd__and2_1
X_4395_ _4401_/A vssd1 vssd1 vccd1 vccd1 _4400_/A sky130_fd_sc_hd__buf_2
XFILLER_58_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6134_ _6134_/A _6134_/B _5941_/X vssd1 vssd1 vccd1 vccd1 _6321_/A sky130_fd_sc_hd__or3b_1
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6065_ _6119_/A vssd1 vssd1 vccd1 vccd1 _6316_/B sky130_fd_sc_hd__clkbuf_2
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5016_ _5016_/A _5120_/A _5126_/B _5044_/C vssd1 vssd1 vccd1 vccd1 _5153_/B sky130_fd_sc_hd__or4_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6967_ _6967_/A _6967_/B _6967_/C vssd1 vssd1 vccd1 vccd1 _7347_/A sky130_fd_sc_hd__and3_1
XFILLER_81_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8706_ _8734_/CLK _8706_/D vssd1 vssd1 vccd1 vccd1 _8706_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5918_ _5919_/A _5919_/B vssd1 vssd1 vccd1 vccd1 _5964_/A sky130_fd_sc_hd__nor2_2
XFILLER_41_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6898_ _6951_/A _6898_/B vssd1 vssd1 vccd1 vccd1 _6952_/B sky130_fd_sc_hd__xnor2_2
X_8637_ _8710_/CLK _8637_/D vssd1 vssd1 vccd1 vccd1 _8637_/Q sky130_fd_sc_hd__dfxtp_1
X_5849_ _5851_/A _5851_/B vssd1 vssd1 vccd1 vccd1 _6060_/A sky130_fd_sc_hd__and2_1
XFILLER_21_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8568_ _8568_/A vssd1 vssd1 vccd1 vccd1 _8733_/D sky130_fd_sc_hd__clkbuf_1
X_7519_ _7520_/A _7526_/B vssd1 vssd1 vccd1 vccd1 _7521_/A sky130_fd_sc_hd__and2_1
X_8499_ _8499_/A _8499_/B vssd1 vssd1 vccd1 vccd1 _8501_/A sky130_fd_sc_hd__xor2_1
XFILLER_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7870_ _8321_/A _8330_/A vssd1 vssd1 vccd1 vccd1 _7880_/A sky130_fd_sc_hd__nor2_1
X_6821_ _7146_/A _7434_/B vssd1 vssd1 vccd1 vccd1 _7095_/A sky130_fd_sc_hd__xor2_1
XFILLER_63_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6752_ _7060_/B vssd1 vssd1 vccd1 vccd1 _7063_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_50_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6683_ _6699_/A _6700_/A _6702_/B _6682_/X vssd1 vssd1 vccd1 vccd1 _6793_/C sky130_fd_sc_hd__a31o_2
X_5703_ _5701_/X _5572_/B _5702_/X vssd1 vssd1 vccd1 vccd1 _5775_/A sky130_fd_sc_hd__a21o_1
XFILLER_31_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8422_ _8422_/A _8422_/B vssd1 vssd1 vccd1 vccd1 _8487_/B sky130_fd_sc_hd__xor2_1
X_5634_ _5634_/A _5634_/B vssd1 vssd1 vccd1 vccd1 _5634_/X sky130_fd_sc_hd__and2_1
X_8353_ _8353_/A _8356_/B vssd1 vssd1 vccd1 vccd1 _8431_/B sky130_fd_sc_hd__xnor2_1
X_7304_ _7304_/A _7304_/B vssd1 vssd1 vccd1 vccd1 _7304_/Y sky130_fd_sc_hd__nor2_1
X_5565_ _5702_/A _5702_/B vssd1 vssd1 vccd1 vccd1 _5572_/A sky130_fd_sc_hd__xnor2_1
X_4516_ _5079_/A _5226_/A vssd1 vssd1 vccd1 vccd1 _4986_/A sky130_fd_sc_hd__or2_1
X_8284_ _8284_/A _8367_/A vssd1 vssd1 vccd1 vccd1 _8291_/B sky130_fd_sc_hd__xnor2_1
XFILLER_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5496_ _5506_/B vssd1 vssd1 vccd1 vccd1 _5780_/C sky130_fd_sc_hd__clkbuf_2
X_4447_ _4449_/A vssd1 vssd1 vccd1 vccd1 _4447_/Y sky130_fd_sc_hd__inv_2
X_7235_ _7235_/A _7235_/B vssd1 vssd1 vccd1 vccd1 _7238_/A sky130_fd_sc_hd__xnor2_1
XFILLER_104_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7166_ _7069_/A _7211_/A _7068_/X vssd1 vssd1 vccd1 vccd1 _7167_/B sky130_fd_sc_hd__o21ba_1
X_4378_ _4382_/A vssd1 vssd1 vccd1 vccd1 _4378_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6117_ _6117_/A _6117_/B vssd1 vssd1 vccd1 vccd1 _6129_/A sky130_fd_sc_hd__nand2_1
X_7097_ _7097_/A _7097_/B vssd1 vssd1 vccd1 vccd1 _7112_/B sky130_fd_sc_hd__xor2_1
XFILLER_58_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6048_ _6048_/A _6052_/B vssd1 vssd1 vccd1 vccd1 _6085_/A sky130_fd_sc_hd__xnor2_1
XFILLER_37_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_8_0_wb_clk_i clkbuf_4_9_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _8695_/CLK
+ sky130_fd_sc_hd__clkbuf_2
X_7999_ _8079_/A _8079_/B vssd1 vssd1 vccd1 vccd1 _8084_/A sky130_fd_sc_hd__xnor2_1
XFILLER_26_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8808__75 vssd1 vssd1 vccd1 vccd1 _8808__75/HI _8917_/A sky130_fd_sc_hd__conb_1
XFILLER_94_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5350_ _5350_/A _5350_/B vssd1 vssd1 vccd1 vccd1 _8649_/D sky130_fd_sc_hd__nor2_1
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5281_ _8631_/Q _5285_/B vssd1 vssd1 vccd1 vccd1 _5281_/X sky130_fd_sc_hd__or2_1
X_7020_ _6902_/A _6950_/X _7018_/Y _7019_/X vssd1 vssd1 vccd1 vccd1 _7302_/A sky130_fd_sc_hd__a211oi_1
XFILLER_4_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7922_ _7922_/A _7922_/B vssd1 vssd1 vccd1 vccd1 _7926_/A sky130_fd_sc_hd__xnor2_1
XFILLER_63_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7853_ _7795_/A _7853_/B vssd1 vssd1 vccd1 vccd1 _7945_/A sky130_fd_sc_hd__and2b_1
X_6804_ _6804_/A _6804_/B _6804_/C vssd1 vssd1 vccd1 vccd1 _6804_/X sky130_fd_sc_hd__and3_1
X_4996_ _4996_/A vssd1 vssd1 vccd1 vccd1 _5016_/A sky130_fd_sc_hd__clkbuf_2
X_7784_ _8228_/A vssd1 vssd1 vccd1 vccd1 _8335_/A sky130_fd_sc_hd__clkbuf_2
X_6735_ _6735_/A _6870_/A _6870_/B vssd1 vssd1 vccd1 vccd1 _7080_/A sky130_fd_sc_hd__and3_1
XFILLER_23_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6666_ _6677_/A _6677_/B vssd1 vssd1 vccd1 vccd1 _6734_/B sky130_fd_sc_hd__xor2_2
X_6597_ _6607_/A _6597_/B vssd1 vssd1 vccd1 vccd1 _6730_/A sky130_fd_sc_hd__nor2_2
X_5617_ _5813_/A _5627_/A vssd1 vssd1 vccd1 vccd1 _6039_/A sky130_fd_sc_hd__nand2_1
X_8405_ _8405_/A _8405_/B vssd1 vssd1 vccd1 vccd1 _8407_/A sky130_fd_sc_hd__nand2_1
X_5548_ _5548_/A _5548_/B _5548_/C vssd1 vssd1 vccd1 vccd1 _5549_/B sky130_fd_sc_hd__nor3_1
X_8336_ _8131_/B _8411_/S _8335_/Y _8221_/A vssd1 vssd1 vccd1 vccd1 _8337_/B sky130_fd_sc_hd__o2bb2a_1
X_8267_ _8269_/A _8269_/B vssd1 vssd1 vccd1 vccd1 _8509_/A sky130_fd_sc_hd__xnor2_1
X_7218_ _7209_/X _7216_/Y _7217_/X _7188_/Y vssd1 vssd1 vccd1 vccd1 _7223_/A sky130_fd_sc_hd__a211oi_1
X_5479_ _5566_/A _5998_/A vssd1 vssd1 vccd1 vccd1 _5479_/Y sky130_fd_sc_hd__nand2_1
X_8198_ _8390_/A _8303_/B vssd1 vssd1 vccd1 vccd1 _8199_/B sky130_fd_sc_hd__xnor2_1
XFILLER_48_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7149_ _7177_/A _7177_/B vssd1 vssd1 vccd1 vccd1 _7157_/A sky130_fd_sc_hd__nand2_1
XFILLER_100_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4850_ _4879_/A _4904_/A _4977_/A vssd1 vssd1 vccd1 vccd1 _5007_/A sky130_fd_sc_hd__o21bai_4
XFILLER_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6520_ _6521_/A _6526_/B vssd1 vssd1 vccd1 vccd1 _6520_/Y sky130_fd_sc_hd__nor2_1
X_4781_ _4781_/A _4781_/B vssd1 vssd1 vccd1 vccd1 _4781_/X sky130_fd_sc_hd__and2_1
XFILLER_20_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6451_ _8690_/Q _6450_/B _6406_/B vssd1 vssd1 vccd1 vccd1 _6452_/B sky130_fd_sc_hd__o21ai_1
X_6382_ _8677_/Q _8678_/Q _8681_/Q _6394_/D vssd1 vssd1 vccd1 vccd1 _6382_/X sky130_fd_sc_hd__o211a_1
X_5402_ _8657_/Q _5402_/B vssd1 vssd1 vccd1 vccd1 _5402_/Y sky130_fd_sc_hd__xnor2_1
X_5333_ _8644_/Q _5332_/B _5323_/X vssd1 vssd1 vccd1 vccd1 _5334_/B sky130_fd_sc_hd__o21ai_1
X_8121_ _8321_/B _8028_/X _8027_/Y _7887_/B vssd1 vssd1 vccd1 vccd1 _8224_/A sky130_fd_sc_hd__a2bb2o_1
X_5264_ _8666_/Q _5258_/X _5263_/X _4651_/X vssd1 vssd1 vccd1 vccd1 _8624_/D sky130_fd_sc_hd__o211a_1
X_8052_ _8052_/A _8368_/B vssd1 vssd1 vccd1 vccd1 _8085_/B sky130_fd_sc_hd__nor2_1
X_7003_ _7003_/A _7003_/B vssd1 vssd1 vccd1 vccd1 _7342_/A sky130_fd_sc_hd__xnor2_1
X_5195_ _5183_/C _5248_/B _5192_/X _5194_/X vssd1 vssd1 vccd1 vccd1 _5195_/X sky130_fd_sc_hd__o31a_1
XFILLER_83_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8799__66 vssd1 vssd1 vccd1 vccd1 _8799__66/HI _8908_/A sky130_fd_sc_hd__conb_1
XFILLER_95_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8885_ _8885_/A _4398_/Y vssd1 vssd1 vccd1 vccd1 io_out[22] sky130_fd_sc_hd__ebufn_8
X_7905_ _8281_/A _7905_/B vssd1 vssd1 vccd1 vccd1 _7919_/A sky130_fd_sc_hd__or2_1
XFILLER_70_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7836_ _7836_/A _8052_/A _7836_/C vssd1 vssd1 vccd1 vccd1 _8514_/A sky130_fd_sc_hd__and3_2
XFILLER_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4979_ _4979_/A _5162_/B vssd1 vssd1 vccd1 vccd1 _4987_/C sky130_fd_sc_hd__or2_1
X_7767_ _7871_/A _8735_/Q vssd1 vssd1 vccd1 vccd1 _7768_/B sky130_fd_sc_hd__and2b_1
X_6718_ _6876_/B _7128_/B _7352_/C vssd1 vssd1 vccd1 vccd1 _6780_/B sky130_fd_sc_hd__or3_1
X_7698_ _7875_/A vssd1 vssd1 vccd1 vccd1 _7885_/A sky130_fd_sc_hd__buf_2
X_6649_ _6797_/A _6980_/A vssd1 vssd1 vccd1 vccd1 _6650_/B sky130_fd_sc_hd__and2_1
X_8319_ _8319_/A _8319_/B vssd1 vssd1 vccd1 vccd1 _8319_/Y sky130_fd_sc_hd__nand2_1
XFILLER_59_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5951_ _5947_/X _6171_/A _5859_/A vssd1 vssd1 vccd1 vccd1 _5953_/B sky130_fd_sc_hd__a21o_1
XFILLER_25_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4902_ _5169_/A _5035_/A vssd1 vssd1 vccd1 vccd1 _5046_/A sky130_fd_sc_hd__or2_1
X_8670_ _8674_/CLK _8670_/D vssd1 vssd1 vccd1 vccd1 _8670_/Q sky130_fd_sc_hd__dfxtp_1
X_5882_ _5881_/B _5882_/B vssd1 vssd1 vccd1 vccd1 _5882_/X sky130_fd_sc_hd__and2b_1
X_4833_ _4878_/A _4904_/B vssd1 vssd1 vccd1 vccd1 _4998_/B sky130_fd_sc_hd__nor2_1
XFILLER_33_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7621_ _8574_/A _7621_/B vssd1 vssd1 vccd1 vccd1 _7621_/Y sky130_fd_sc_hd__nor2_1
X_4764_ _4828_/C _4898_/A vssd1 vssd1 vccd1 vccd1 _4786_/C sky130_fd_sc_hd__nor2_2
X_7552_ _8734_/Q vssd1 vssd1 vccd1 vccd1 _8571_/A sky130_fd_sc_hd__clkbuf_2
X_6503_ _6503_/A _7548_/B vssd1 vssd1 vccd1 vccd1 _6507_/A sky130_fd_sc_hd__nor2_1
X_7483_ _7475_/A _7479_/B _7475_/C _7202_/A vssd1 vssd1 vccd1 vccd1 _7484_/A sky130_fd_sc_hd__a31o_1
X_6434_ _6437_/C _6434_/B vssd1 vssd1 vccd1 vccd1 _8684_/D sky130_fd_sc_hd__nor2_1
X_4695_ _4700_/A _4694_/X _4727_/A vssd1 vssd1 vccd1 vccd1 _8604_/D sky130_fd_sc_hd__a21boi_1
X_6365_ _5398_/A _6363_/Y _6373_/S _5397_/X _6360_/A vssd1 vssd1 vccd1 vccd1 _8672_/D
+ sky130_fd_sc_hd__a32o_1
X_5316_ _5323_/A vssd1 vssd1 vccd1 vccd1 _5362_/A sky130_fd_sc_hd__clkbuf_2
X_6296_ _6299_/B _6296_/B vssd1 vssd1 vccd1 vccd1 _6296_/X sky130_fd_sc_hd__and2_1
X_8104_ _8018_/Y _8503_/B _8506_/B _8506_/A _8506_/C vssd1 vssd1 vccd1 vccd1 _8509_/B
+ sky130_fd_sc_hd__o2111ai_4
X_5247_ _5038_/A _5243_/X _5236_/X _5244_/X _5246_/X vssd1 vssd1 vccd1 vccd1 _5248_/C
+ sky130_fd_sc_hd__o32a_1
X_8035_ _8410_/A vssd1 vssd1 vccd1 vccd1 _8325_/A sky130_fd_sc_hd__buf_2
XFILLER_29_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5178_ _5172_/X _5177_/X _4698_/B _4960_/B vssd1 vssd1 vccd1 vccd1 _5178_/X sky130_fd_sc_hd__a211o_1
XFILLER_28_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8937_ _8937_/A _4459_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[36] sky130_fd_sc_hd__ebufn_8
XFILLER_71_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8868_ _8868_/A _4378_/Y vssd1 vssd1 vccd1 vccd1 io_out[5] sky130_fd_sc_hd__ebufn_8
XFILLER_71_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7819_ _7819_/A _7819_/B vssd1 vssd1 vccd1 vccd1 _7822_/A sky130_fd_sc_hd__xnor2_1
XFILLER_20_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4480_ _4720_/A _4714_/A _4480_/C vssd1 vssd1 vccd1 vccd1 _4718_/A sky130_fd_sc_hd__and3_1
XFILLER_7_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6150_ _6300_/B _6150_/B vssd1 vssd1 vccd1 vccd1 _6311_/B sky130_fd_sc_hd__xnor2_1
X_5101_ _5212_/A _5116_/A _5173_/B vssd1 vssd1 vccd1 vccd1 _5102_/B sky130_fd_sc_hd__or3b_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_10_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8689_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6081_ _6046_/B _6079_/X _6078_/Y _6072_/X vssd1 vssd1 vccd1 vccd1 _6083_/B sky130_fd_sc_hd__o211a_1
X_5032_ _4930_/X _4973_/X _4988_/X _5031_/X vssd1 vssd1 vccd1 vccd1 _5032_/X sky130_fd_sc_hd__a31o_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8769__36 vssd1 vssd1 vccd1 vccd1 _8769__36/HI _8864_/A sky130_fd_sc_hd__conb_1
XFILLER_65_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6983_ _7369_/A _7369_/B vssd1 vssd1 vccd1 vccd1 _6984_/B sky130_fd_sc_hd__xor2_1
XFILLER_25_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5934_ _5926_/A _5926_/B _5933_/Y vssd1 vssd1 vccd1 vccd1 _6161_/B sky130_fd_sc_hd__a21o_1
XFILLER_15_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8722_ _8732_/CLK _8722_/D vssd1 vssd1 vccd1 vccd1 _8722_/Q sky130_fd_sc_hd__dfxtp_1
X_8653_ _8715_/CLK _8653_/D vssd1 vssd1 vccd1 vccd1 _8653_/Q sky130_fd_sc_hd__dfxtp_1
X_5865_ _6196_/A _5866_/B vssd1 vssd1 vccd1 vccd1 _5979_/A sky130_fd_sc_hd__and2_1
X_4816_ _4979_/A _5192_/B vssd1 vssd1 vccd1 vccd1 _5111_/B sky130_fd_sc_hd__or2_1
XFILLER_21_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7604_ _7597_/A _7599_/B _7597_/B vssd1 vssd1 vccd1 vccd1 _7604_/X sky130_fd_sc_hd__o21ba_1
XFILLER_21_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5796_ _5796_/A _5872_/C vssd1 vssd1 vccd1 vccd1 _5798_/B sky130_fd_sc_hd__xnor2_1
X_8584_ _8672_/CLK _8584_/D vssd1 vssd1 vccd1 vccd1 _8584_/Q sky130_fd_sc_hd__dfxtp_1
X_7535_ _7535_/A _7535_/B _7535_/C vssd1 vssd1 vccd1 vccd1 _7547_/S sky130_fd_sc_hd__or3_2
X_4747_ _4828_/C _5263_/B _4740_/B _4900_/A _4746_/X vssd1 vssd1 vccd1 vccd1 _8613_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_31_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7466_ _7466_/A _7466_/B vssd1 vssd1 vccd1 vccd1 _7467_/B sky130_fd_sc_hd__xnor2_2
X_4678_ _4960_/A vssd1 vssd1 vccd1 vccd1 _4702_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6417_ _6394_/D _6418_/C _6416_/Y vssd1 vssd1 vccd1 vccd1 _8679_/D sky130_fd_sc_hd__a21oi_1
X_7397_ _7397_/A _7397_/B vssd1 vssd1 vccd1 vccd1 _7397_/X sky130_fd_sc_hd__or2_1
X_6348_ _6338_/S _6343_/B _6342_/A vssd1 vssd1 vccd1 vccd1 _6350_/B sky130_fd_sc_hd__o21a_1
XFILLER_88_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6279_ _6229_/A _6277_/Y _6278_/Y vssd1 vssd1 vccd1 vccd1 _6280_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8018_ _8503_/A vssd1 vssd1 vccd1 vccd1 _8018_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8783__50 vssd1 vssd1 vccd1 vccd1 _8783__50/HI _8892_/A sky130_fd_sc_hd__conb_1
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5650_ _5746_/B _6097_/B _5687_/A _6049_/A vssd1 vssd1 vccd1 vccd1 _5729_/A sky130_fd_sc_hd__a31o_1
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4601_ _8586_/Q _4604_/C vssd1 vssd1 vccd1 vccd1 _4603_/A sky130_fd_sc_hd__and2_1
X_5581_ _5723_/A _5581_/B vssd1 vssd1 vccd1 vccd1 _5582_/B sky130_fd_sc_hd__xnor2_1
X_7320_ _7403_/A _7320_/B vssd1 vssd1 vccd1 vccd1 _7321_/B sky130_fd_sc_hd__xnor2_1
X_4532_ _4828_/A vssd1 vssd1 vccd1 vccd1 _4758_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4463_ _4464_/A vssd1 vssd1 vccd1 vccd1 _4463_/Y sky130_fd_sc_hd__inv_2
X_7251_ _7249_/A _7248_/C _7248_/B vssd1 vssd1 vccd1 vccd1 _7286_/B sky130_fd_sc_hd__a21o_1
XFILLER_7_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6202_ _6202_/A _6202_/B vssd1 vssd1 vccd1 vccd1 _6202_/X sky130_fd_sc_hd__and2_1
X_7182_ _7182_/A _7182_/B vssd1 vssd1 vccd1 vccd1 _7208_/B sky130_fd_sc_hd__xor2_1
X_4394_ _4394_/A vssd1 vssd1 vccd1 vccd1 _4394_/Y sky130_fd_sc_hd__inv_2
X_6133_ _6133_/A _6133_/B vssd1 vssd1 vccd1 vccd1 _6297_/A sky130_fd_sc_hd__xnor2_1
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6064_ _6033_/X _6096_/B _6036_/B vssd1 vssd1 vccd1 vccd1 _6075_/B sky130_fd_sc_hd__o21ai_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5015_ _5229_/B _5022_/B _5128_/B vssd1 vssd1 vccd1 vccd1 _5015_/X sky130_fd_sc_hd__or3_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6966_ _6880_/X _6879_/A _7443_/B _6882_/B vssd1 vssd1 vccd1 vccd1 _6967_/C sky130_fd_sc_hd__a22o_1
XFILLER_81_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8705_ _8734_/CLK _8705_/D vssd1 vssd1 vccd1 vccd1 _8705_/Q sky130_fd_sc_hd__dfxtp_1
X_5917_ _5841_/A _5840_/B _5838_/Y vssd1 vssd1 vccd1 vccd1 _5919_/B sky130_fd_sc_hd__a21o_1
X_6897_ _6897_/A _6987_/B vssd1 vssd1 vccd1 vccd1 _6898_/B sky130_fd_sc_hd__xnor2_1
XFILLER_42_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8636_ _8710_/CLK _8636_/D vssd1 vssd1 vccd1 vccd1 _8636_/Q sky130_fd_sc_hd__dfxtp_1
X_5848_ _5848_/A _5848_/B vssd1 vssd1 vccd1 vccd1 _5851_/B sky130_fd_sc_hd__xor2_1
X_8567_ _8567_/A _8567_/B vssd1 vssd1 vccd1 vccd1 _8568_/A sky130_fd_sc_hd__and2_1
X_5779_ _5713_/X _5711_/B _5778_/Y vssd1 vssd1 vccd1 vccd1 _5881_/B sky130_fd_sc_hd__a21oi_1
X_7518_ _7514_/A _5362_/X _6508_/X _7517_/X vssd1 vssd1 vccd1 vccd1 _8710_/D sky130_fd_sc_hd__a22o_1
X_8498_ _8495_/Y _8496_/X _8497_/X vssd1 vssd1 vccd1 vccd1 _8512_/C sky130_fd_sc_hd__o21ai_1
X_7449_ _7449_/A _7449_/B vssd1 vssd1 vccd1 vccd1 _7450_/B sky130_fd_sc_hd__nand2_1
XFILLER_89_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6820_ _6865_/B _6820_/B vssd1 vssd1 vccd1 vccd1 _7115_/A sky130_fd_sc_hd__xnor2_1
XFILLER_50_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6751_ _7335_/B _7173_/A vssd1 vssd1 vccd1 vccd1 _6856_/A sky130_fd_sc_hd__nand2_1
Xclkbuf_1_1_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
X_6682_ _6715_/A _7172_/B _7130_/A vssd1 vssd1 vccd1 vccd1 _6682_/X sky130_fd_sc_hd__and3_1
X_5702_ _5702_/A _5702_/B vssd1 vssd1 vccd1 vccd1 _5702_/X sky130_fd_sc_hd__and2_1
X_8421_ _8421_/A _8421_/B vssd1 vssd1 vccd1 vccd1 _8422_/B sky130_fd_sc_hd__xnor2_1
X_5633_ _5746_/B _5859_/B vssd1 vssd1 vccd1 vccd1 _5685_/A sky130_fd_sc_hd__nand2_1
XFILLER_31_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8352_ _8355_/B _8352_/B vssd1 vssd1 vccd1 vccd1 _8356_/B sky130_fd_sc_hd__xnor2_1
X_5564_ _5893_/B _5564_/B vssd1 vssd1 vccd1 vccd1 _5702_/B sky130_fd_sc_hd__xnor2_1
X_7303_ _7303_/A vssd1 vssd1 vccd1 vccd1 _7303_/Y sky130_fd_sc_hd__inv_2
X_4515_ _8604_/Q vssd1 vssd1 vccd1 vccd1 _5226_/A sky130_fd_sc_hd__clkbuf_2
X_8283_ _8283_/A vssd1 vssd1 vccd1 vccd1 _8367_/A sky130_fd_sc_hd__buf_2
X_5495_ _5493_/A _5493_/C _5493_/B vssd1 vssd1 vccd1 vccd1 _5506_/B sky130_fd_sc_hd__a21o_1
X_4446_ _4449_/A vssd1 vssd1 vccd1 vccd1 _4446_/Y sky130_fd_sc_hd__inv_2
X_7234_ _7234_/A _7234_/B vssd1 vssd1 vccd1 vccd1 _7235_/A sky130_fd_sc_hd__nor2_1
X_4377_ _4401_/A vssd1 vssd1 vccd1 vccd1 _4382_/A sky130_fd_sc_hd__clkbuf_4
X_7165_ _7173_/A _7165_/B vssd1 vssd1 vccd1 vccd1 _7212_/A sky130_fd_sc_hd__xnor2_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6116_ _6116_/A _6116_/B vssd1 vssd1 vccd1 vccd1 _6117_/B sky130_fd_sc_hd__nand2_1
XFILLER_85_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7096_ _7096_/A _7096_/B vssd1 vssd1 vccd1 vccd1 _7097_/B sky130_fd_sc_hd__and2_1
XFILLER_58_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6047_ _6047_/A _6047_/B vssd1 vssd1 vccd1 vccd1 _6052_/B sky130_fd_sc_hd__xor2_1
XFILLER_39_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7998_ _7998_/A _7998_/B vssd1 vssd1 vccd1 vccd1 _8079_/B sky130_fd_sc_hd__xnor2_1
XFILLER_41_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8753__20 vssd1 vssd1 vccd1 vccd1 _8753__20/HI _8848_/A sky130_fd_sc_hd__conb_1
X_6949_ _6949_/A _6949_/B vssd1 vssd1 vccd1 vccd1 _6949_/Y sky130_fd_sc_hd__nor2_1
XFILLER_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8619_ _8733_/CLK _8619_/D vssd1 vssd1 vccd1 vccd1 _8619_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5280_ _8705_/Q _5271_/X _5278_/X _5279_/X vssd1 vssd1 vccd1 vccd1 _8630_/D sky130_fd_sc_hd__o211a_1
XFILLER_4_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7921_ _7985_/B _7921_/B vssd1 vssd1 vccd1 vccd1 _7922_/B sky130_fd_sc_hd__xnor2_1
XFILLER_82_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7852_ _7852_/A vssd1 vssd1 vccd1 vccd1 _7852_/Y sky130_fd_sc_hd__inv_2
X_4995_ _5120_/A vssd1 vssd1 vccd1 vccd1 _5215_/B sky130_fd_sc_hd__clkbuf_2
X_6803_ _6804_/C _6803_/B vssd1 vssd1 vccd1 vccd1 _6803_/X sky130_fd_sc_hd__and2b_1
X_7783_ _7783_/A vssd1 vssd1 vccd1 vccd1 _8228_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6734_ _6734_/A _6734_/B vssd1 vssd1 vccd1 vccd1 _7133_/A sky130_fd_sc_hd__nor2_2
XFILLER_51_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6665_ _6659_/A _6652_/B _6635_/B _6664_/X vssd1 vssd1 vccd1 vccd1 _6677_/B sky130_fd_sc_hd__a31o_1
X_8404_ _8404_/A _8404_/B _8404_/C vssd1 vssd1 vccd1 vccd1 _8405_/B sky130_fd_sc_hd__or3_1
X_6596_ _7548_/A _6596_/B vssd1 vssd1 vccd1 vccd1 _6597_/B sky130_fd_sc_hd__nor2_1
X_5616_ _5642_/A _5642_/B vssd1 vssd1 vccd1 vccd1 _5627_/A sky130_fd_sc_hd__nand2_1
X_5547_ _5548_/A _5548_/B _5548_/C vssd1 vssd1 vccd1 vccd1 _5584_/A sky130_fd_sc_hd__o21a_2
X_8335_ _8335_/A _8410_/B vssd1 vssd1 vccd1 vccd1 _8335_/Y sky130_fd_sc_hd__nor2_1
X_8266_ _8266_/A _8266_/B vssd1 vssd1 vccd1 vccd1 _8269_/B sky130_fd_sc_hd__xnor2_1
X_5478_ _5481_/B vssd1 vssd1 vccd1 vccd1 _5998_/A sky130_fd_sc_hd__clkbuf_2
X_4429_ _4431_/A vssd1 vssd1 vccd1 vccd1 _4429_/Y sky130_fd_sc_hd__clkinv_4
X_7217_ _7188_/A _7188_/B _7188_/C vssd1 vssd1 vccd1 vccd1 _7217_/X sky130_fd_sc_hd__o21a_1
XFILLER_59_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8197_ _8473_/S _8196_/X _8147_/X vssd1 vssd1 vccd1 vccd1 _8303_/B sky130_fd_sc_hd__a21o_1
XFILLER_86_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7148_ _7148_/A _7148_/B vssd1 vssd1 vccd1 vccd1 _7177_/B sky130_fd_sc_hd__nor2_1
XFILLER_48_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7079_ _7145_/B _7138_/B _7078_/Y vssd1 vssd1 vccd1 vccd1 _7105_/A sky130_fd_sc_hd__a21o_1
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4780_ _4781_/A _4781_/B _4779_/Y _4651_/X vssd1 vssd1 vccd1 vccd1 _8619_/D sky130_fd_sc_hd__o211a_1
XFILLER_33_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6450_ _8690_/Q _6450_/B vssd1 vssd1 vccd1 vccd1 _6455_/C sky130_fd_sc_hd__and2_1
X_6381_ _8679_/Q vssd1 vssd1 vccd1 vccd1 _6394_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_5401_ _5401_/A _5401_/B vssd1 vssd1 vccd1 vccd1 _5402_/B sky130_fd_sc_hd__nand2_1
X_5332_ _8644_/Q _5332_/B vssd1 vssd1 vccd1 vccd1 _5338_/C sky130_fd_sc_hd__and2_1
X_8120_ _8203_/B _8120_/B vssd1 vssd1 vccd1 vccd1 _8126_/A sky130_fd_sc_hd__xnor2_1
XFILLER_102_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5263_ _8624_/Q _5263_/B vssd1 vssd1 vccd1 vccd1 _5263_/X sky130_fd_sc_hd__or2_1
X_8051_ _8051_/A _8071_/A vssd1 vssd1 vccd1 vccd1 _8368_/B sky130_fd_sc_hd__nand2_1
X_7002_ _7002_/A _7329_/B vssd1 vssd1 vccd1 vccd1 _7003_/B sky130_fd_sc_hd__xor2_1
X_5194_ _5194_/A _5209_/B _5194_/C _5208_/C vssd1 vssd1 vccd1 vccd1 _5194_/X sky130_fd_sc_hd__or4_1
XFILLER_68_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8884_ _8884_/A _4397_/Y vssd1 vssd1 vccd1 vccd1 io_out[21] sky130_fd_sc_hd__ebufn_8
XFILLER_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7904_ _7813_/B _7809_/B _7903_/X vssd1 vssd1 vccd1 vccd1 _7914_/A sky130_fd_sc_hd__a21oi_1
XFILLER_24_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7835_ _7835_/A _7835_/B vssd1 vssd1 vccd1 vccd1 _7836_/C sky130_fd_sc_hd__nand2_1
XFILLER_24_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4978_ _5185_/B _5190_/B _5107_/A vssd1 vssd1 vccd1 vccd1 _5162_/B sky130_fd_sc_hd__or3_1
XFILLER_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7766_ _8735_/Q _7871_/A vssd1 vssd1 vccd1 vccd1 _7768_/A sky130_fd_sc_hd__and2b_1
X_6717_ _6972_/C vssd1 vssd1 vccd1 vccd1 _7128_/B sky130_fd_sc_hd__clkbuf_2
X_7697_ _8118_/A _7728_/A vssd1 vssd1 vccd1 vccd1 _7875_/A sky130_fd_sc_hd__nand2_1
X_6648_ _6797_/A _6980_/A vssd1 vssd1 vccd1 vccd1 _6768_/A sky130_fd_sc_hd__nor2_1
X_6579_ _6579_/A _6579_/B vssd1 vssd1 vccd1 vccd1 _6670_/A sky130_fd_sc_hd__xnor2_1
XFILLER_3_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8318_ _8237_/A _8345_/B _8236_/B _8238_/B _8238_/A vssd1 vssd1 vccd1 vccd1 _8384_/A
+ sky130_fd_sc_hd__a32oi_4
XFILLER_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8249_ _8277_/A _8277_/B vssd1 vssd1 vccd1 vccd1 _8250_/B sky130_fd_sc_hd__xor2_1
XFILLER_59_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5950_ _5953_/A _6119_/B vssd1 vssd1 vccd1 vccd1 _6171_/A sky130_fd_sc_hd__nand2_1
X_4901_ _5193_/A _5238_/C vssd1 vssd1 vccd1 vccd1 _5035_/A sky130_fd_sc_hd__or2_1
XFILLER_33_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5881_ _5882_/B _5881_/B vssd1 vssd1 vccd1 vccd1 _5881_/X sky130_fd_sc_hd__and2b_1
X_7620_ _7620_/A _7620_/B vssd1 vssd1 vccd1 vccd1 _7621_/B sky130_fd_sc_hd__xnor2_1
X_4832_ _5223_/B _5044_/B vssd1 vssd1 vccd1 vccd1 _4966_/A sky130_fd_sc_hd__or2_1
X_7551_ _7551_/A vssd1 vssd1 vccd1 vccd1 _8715_/D sky130_fd_sc_hd__clkbuf_1
X_4763_ _4763_/A _4763_/B vssd1 vssd1 vccd1 vccd1 _4765_/B sky130_fd_sc_hd__nand2_1
XFILLER_21_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6502_ _6502_/A vssd1 vssd1 vccd1 vccd1 _7548_/B sky130_fd_sc_hd__clkbuf_2
X_4694_ _4694_/A _4711_/A vssd1 vssd1 vccd1 vccd1 _4694_/X sky130_fd_sc_hd__or2_1
X_7482_ _7482_/A _7482_/B vssd1 vssd1 vccd1 vccd1 _7482_/Y sky130_fd_sc_hd__nand2_1
X_6433_ _8684_/Q _6431_/A _6406_/B vssd1 vssd1 vccd1 vccd1 _6434_/B sky130_fd_sc_hd__o21ai_1
X_6364_ _6364_/A _6364_/B vssd1 vssd1 vccd1 vccd1 _6373_/S sky130_fd_sc_hd__or2_1
X_5315_ _8637_/Q _6466_/B _5307_/B _8639_/Q vssd1 vssd1 vccd1 vccd1 _5317_/B sky130_fd_sc_hd__a31o_1
X_6295_ _6295_/A _6298_/A vssd1 vssd1 vccd1 vccd1 _6296_/B sky130_fd_sc_hd__nand2_1
X_8103_ _8101_/A _8102_/B _8503_/A _8100_/X vssd1 vssd1 vccd1 vccd1 _8506_/C sky130_fd_sc_hd__a2bb2o_1
XFILLER_102_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5246_ _5233_/B _5007_/B _5179_/X _5245_/X _5038_/A vssd1 vssd1 vccd1 vccd1 _5246_/X
+ sky130_fd_sc_hd__o32a_1
X_8034_ _8034_/A vssd1 vssd1 vccd1 vccd1 _8321_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_29_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5177_ _5212_/A _5202_/C _5177_/C vssd1 vssd1 vccd1 vccd1 _5177_/X sky130_fd_sc_hd__or3_1
X_8936_ _8936_/A _4458_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[35] sky130_fd_sc_hd__ebufn_8
XFILLER_83_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8867_ _8867_/A _4375_/Y vssd1 vssd1 vccd1 vccd1 io_out[4] sky130_fd_sc_hd__ebufn_8
XFILLER_101_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7818_ _7818_/A _7818_/B vssd1 vssd1 vccd1 vccd1 _7819_/B sky130_fd_sc_hd__xnor2_1
X_7749_ _7675_/A _7675_/B _7748_/Y _7661_/X vssd1 vssd1 vccd1 vccd1 _7850_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_94_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6080_ _6072_/X _6078_/Y _6079_/X _6046_/B vssd1 vssd1 vccd1 vccd1 _6084_/A sky130_fd_sc_hd__a211oi_2
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5100_ _5100_/A _5100_/B vssd1 vssd1 vccd1 vccd1 _5116_/A sky130_fd_sc_hd__nand2_1
XFILLER_97_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5031_ _5056_/A _5024_/X _5028_/X _5096_/A vssd1 vssd1 vccd1 vccd1 _5031_/X sky130_fd_sc_hd__o211a_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6982_ _7031_/S vssd1 vssd1 vccd1 vccd1 _7369_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_80_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8721_ _8732_/CLK _8721_/D vssd1 vssd1 vccd1 vccd1 _8721_/Q sky130_fd_sc_hd__dfxtp_1
X_5933_ _5933_/A _5933_/B vssd1 vssd1 vccd1 vccd1 _5933_/Y sky130_fd_sc_hd__nor2_1
X_8652_ _8677_/CLK _8652_/D vssd1 vssd1 vccd1 vccd1 _8652_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5864_ _6194_/A _5862_/Y _5863_/Y vssd1 vssd1 vccd1 vccd1 _5866_/B sky130_fd_sc_hd__a21oi_1
XFILLER_33_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4815_ _4919_/A _4827_/A vssd1 vssd1 vccd1 vccd1 _5192_/B sky130_fd_sc_hd__nor2_1
XFILLER_33_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7603_ _8721_/Q _7617_/B vssd1 vssd1 vccd1 vccd1 _7603_/X sky130_fd_sc_hd__xor2_1
X_8583_ _8672_/CLK _8583_/D vssd1 vssd1 vccd1 vccd1 _8583_/Q sky130_fd_sc_hd__dfxtp_1
X_7534_ _7527_/B _7534_/B vssd1 vssd1 vccd1 vccd1 _7535_/C sky130_fd_sc_hd__and2b_1
X_5795_ _5795_/A _5795_/B vssd1 vssd1 vccd1 vccd1 _5872_/C sky130_fd_sc_hd__xor2_1
X_4746_ _8567_/A vssd1 vssd1 vccd1 vccd1 _4746_/X sky130_fd_sc_hd__clkbuf_4
X_7465_ _7465_/A _7465_/B vssd1 vssd1 vccd1 vccd1 _7466_/B sky130_fd_sc_hd__xnor2_1
X_4677_ _5143_/A vssd1 vssd1 vccd1 vccd1 _4960_/A sky130_fd_sc_hd__clkbuf_2
X_6416_ _6394_/D _6418_/C _6401_/B vssd1 vssd1 vccd1 vccd1 _6416_/Y sky130_fd_sc_hd__o21ai_1
X_7396_ _7397_/A _7397_/B _7395_/X vssd1 vssd1 vccd1 vccd1 _7396_/X sky130_fd_sc_hd__a21bo_1
X_6347_ _6355_/A _6347_/B vssd1 vssd1 vccd1 vccd1 _6350_/A sky130_fd_sc_hd__nand2_1
XFILLER_88_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6278_ _6278_/A _6278_/B vssd1 vssd1 vccd1 vccd1 _6278_/Y sky130_fd_sc_hd__nand2_1
X_5229_ _5229_/A _5229_/B _5229_/C _5229_/D vssd1 vssd1 vccd1 vccd1 _5229_/X sky130_fd_sc_hd__or4_1
XFILLER_69_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8017_ _8017_/A _8017_/B _8017_/C vssd1 vssd1 vccd1 vccd1 _8503_/A sky130_fd_sc_hd__nand3_2
XFILLER_84_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8919_ _8919_/A _4437_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[18] sky130_fd_sc_hd__ebufn_8
XFILLER_71_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_2_3_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_79_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4600_ _4604_/C _4600_/B vssd1 vssd1 vccd1 vccd1 _8585_/D sky130_fd_sc_hd__nor2_1
X_5580_ _5580_/A _5722_/A vssd1 vssd1 vccd1 vccd1 _5581_/B sky130_fd_sc_hd__xnor2_1
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4531_ _4839_/A vssd1 vssd1 vccd1 vccd1 _4828_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4462_ _4464_/A vssd1 vssd1 vccd1 vccd1 _4462_/Y sky130_fd_sc_hd__inv_2
X_7250_ _7250_/A _7289_/A vssd1 vssd1 vccd1 vccd1 _7481_/A sky130_fd_sc_hd__xor2_1
XFILLER_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6201_ _6201_/A _6201_/B vssd1 vssd1 vccd1 vccd1 _6278_/A sky130_fd_sc_hd__nand2_2
XFILLER_98_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8829__96 vssd1 vssd1 vccd1 vccd1 _8829__96/HI _8938_/A sky130_fd_sc_hd__conb_1
X_7181_ _7181_/A _7181_/B vssd1 vssd1 vccd1 vccd1 _7208_/A sky130_fd_sc_hd__xor2_1
X_4393_ _4394_/A vssd1 vssd1 vccd1 vccd1 _4393_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6132_ _6146_/A _6146_/B vssd1 vssd1 vccd1 vccd1 _6295_/A sky130_fd_sc_hd__xnor2_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6063_ _6063_/A _6063_/B vssd1 vssd1 vccd1 vccd1 _6075_/A sky130_fd_sc_hd__xnor2_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5014_ _4891_/C _4948_/B _4937_/A vssd1 vssd1 vccd1 vccd1 _5128_/B sky130_fd_sc_hd__a21oi_4
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6965_ _6964_/B _6964_/C _6964_/A vssd1 vssd1 vccd1 vccd1 _6967_/B sky130_fd_sc_hd__a21o_1
XFILLER_26_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8704_ _8714_/CLK _8704_/D vssd1 vssd1 vccd1 vccd1 _8704_/Q sky130_fd_sc_hd__dfxtp_1
X_5916_ _5937_/A _5916_/B vssd1 vssd1 vccd1 vccd1 _5919_/A sky130_fd_sc_hd__xor2_1
X_6896_ _6954_/A _7327_/A vssd1 vssd1 vccd1 vccd1 _6987_/B sky130_fd_sc_hd__xor2_1
X_8635_ _8715_/CLK _8635_/D vssd1 vssd1 vccd1 vccd1 _8635_/Q sky130_fd_sc_hd__dfxtp_1
X_5847_ _5847_/A _5847_/B vssd1 vssd1 vccd1 vccd1 _5848_/B sky130_fd_sc_hd__xor2_1
XFILLER_21_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8566_ _8565_/X _8576_/A _8566_/S vssd1 vssd1 vccd1 vccd1 _8567_/B sky130_fd_sc_hd__mux2_1
X_5778_ _5778_/A _5802_/A vssd1 vssd1 vccd1 vccd1 _5778_/Y sky130_fd_sc_hd__nor2_1
X_7517_ _7515_/Y _7517_/B vssd1 vssd1 vccd1 vccd1 _7517_/X sky130_fd_sc_hd__and2b_1
X_4729_ _4733_/S _4730_/B vssd1 vssd1 vccd1 vccd1 _4729_/X sky130_fd_sc_hd__and2_1
X_8497_ _8497_/A _8497_/B vssd1 vssd1 vccd1 vccd1 _8497_/X sky130_fd_sc_hd__xor2_1
X_7448_ _7455_/B _7447_/B _7447_/C _7447_/D vssd1 vssd1 vccd1 vccd1 _7449_/B sky130_fd_sc_hd__a22o_1
X_7379_ _7378_/A _7378_/B _7378_/C _7378_/D vssd1 vssd1 vccd1 vccd1 _7379_/X sky130_fd_sc_hd__o22a_1
XFILLER_76_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6750_ _7065_/A _7332_/B vssd1 vssd1 vccd1 vccd1 _7173_/A sky130_fd_sc_hd__nor2_4
XFILLER_63_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5701_ _5702_/A _5702_/B vssd1 vssd1 vccd1 vccd1 _5701_/X sky130_fd_sc_hd__or2_1
X_6681_ _6957_/B vssd1 vssd1 vccd1 vccd1 _7172_/B sky130_fd_sc_hd__clkbuf_2
X_8420_ _8481_/A _8420_/B vssd1 vssd1 vccd1 vccd1 _8421_/B sky130_fd_sc_hd__xnor2_1
X_5632_ _5948_/A vssd1 vssd1 vccd1 vccd1 _5859_/B sky130_fd_sc_hd__clkbuf_2
X_8351_ _8351_/A _8351_/B vssd1 vssd1 vccd1 vccd1 _8352_/B sky130_fd_sc_hd__xnor2_1
X_5563_ _5892_/A _5896_/A _5571_/A _5578_/A vssd1 vssd1 vccd1 vccd1 _5564_/B sky130_fd_sc_hd__o22a_1
X_7302_ _7302_/A _7042_/X vssd1 vssd1 vccd1 vccd1 _7463_/A sky130_fd_sc_hd__or2b_1
X_4514_ _7695_/B vssd1 vssd1 vccd1 vccd1 _5079_/A sky130_fd_sc_hd__clkbuf_2
X_8282_ _8281_/Y _8514_/A _8166_/X vssd1 vssd1 vccd1 vccd1 _8290_/A sky130_fd_sc_hd__o21ai_1
X_5494_ _5506_/A vssd1 vssd1 vccd1 vccd1 _5780_/B sky130_fd_sc_hd__clkbuf_2
X_4445_ _4449_/A vssd1 vssd1 vccd1 vccd1 _4445_/Y sky130_fd_sc_hd__inv_2
X_7233_ _7233_/A _7233_/B vssd1 vssd1 vccd1 vccd1 _7252_/B sky130_fd_sc_hd__xnor2_1
X_4376_ input1/X vssd1 vssd1 vccd1 vccd1 _4401_/A sky130_fd_sc_hd__buf_2
X_7164_ _7293_/A _7292_/B vssd1 vssd1 vccd1 vccd1 _7201_/A sky130_fd_sc_hd__xnor2_1
XFILLER_58_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6115_ _6143_/B _6115_/B vssd1 vssd1 vccd1 vccd1 _6146_/A sky130_fd_sc_hd__and2_1
X_7095_ _7095_/A _7095_/B vssd1 vssd1 vccd1 vccd1 _7096_/B sky130_fd_sc_hd__or2_1
XFILLER_58_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6046_ _6046_/A _6046_/B vssd1 vssd1 vccd1 vccd1 _6048_/A sky130_fd_sc_hd__nor2_1
XFILLER_37_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8742__9 vssd1 vssd1 vccd1 vccd1 _8742__9/HI _8837_/A sky130_fd_sc_hd__conb_1
X_7997_ _8072_/A _8308_/A vssd1 vssd1 vccd1 vccd1 _7998_/B sky130_fd_sc_hd__or2_1
X_6948_ _6948_/A _6948_/B vssd1 vssd1 vccd1 vccd1 _6948_/X sky130_fd_sc_hd__and2_1
XFILLER_53_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6879_ _6879_/A vssd1 vssd1 vccd1 vccd1 _6879_/Y sky130_fd_sc_hd__inv_2
X_8618_ _8733_/CLK _8618_/D vssd1 vssd1 vccd1 vccd1 _8618_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8549_ _7695_/A _8542_/B _8541_/A vssd1 vssd1 vccd1 vccd1 _8550_/B sky130_fd_sc_hd__o21ai_1
XFILLER_1_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7920_ _8008_/B _7920_/B vssd1 vssd1 vccd1 vccd1 _7921_/B sky130_fd_sc_hd__nor2_1
X_7851_ _7851_/A _7851_/B vssd1 vssd1 vccd1 vccd1 _7851_/X sky130_fd_sc_hd__or2_1
X_6802_ _6802_/A _6802_/B vssd1 vssd1 vccd1 vccd1 _6806_/A sky130_fd_sc_hd__xor2_1
XFILLER_63_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4994_ _5227_/A vssd1 vssd1 vccd1 vccd1 _5120_/A sky130_fd_sc_hd__clkbuf_2
X_7782_ _7785_/A _8118_/B _8118_/C vssd1 vssd1 vccd1 vccd1 _7783_/A sky130_fd_sc_hd__and3_1
X_6733_ _7060_/A _7054_/B vssd1 vssd1 vccd1 vccd1 _7091_/A sky130_fd_sc_hd__nor2_1
X_6664_ _6531_/A _7652_/B vssd1 vssd1 vccd1 vccd1 _6664_/X sky130_fd_sc_hd__and2b_1
X_8403_ _8404_/A _8404_/B _8404_/C vssd1 vssd1 vccd1 vccd1 _8405_/A sky130_fd_sc_hd__o21ai_1
X_5615_ _5615_/A _7630_/B vssd1 vssd1 vccd1 vccd1 _5642_/B sky130_fd_sc_hd__nand2_1
X_6595_ _7548_/A _6596_/B vssd1 vssd1 vccd1 vccd1 _6607_/A sky130_fd_sc_hd__and2_1
XFILLER_3_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5546_ _5575_/A _5574_/A _5545_/Y vssd1 vssd1 vccd1 vccd1 _5548_/C sky130_fd_sc_hd__a21oi_1
X_8334_ _8338_/A vssd1 vssd1 vccd1 vccd1 _8411_/S sky130_fd_sc_hd__dlymetal6s2s_1
X_8265_ _8265_/A _8265_/B vssd1 vssd1 vccd1 vccd1 _8269_/A sky130_fd_sc_hd__nand2_1
X_5477_ _5477_/A _5477_/B vssd1 vssd1 vccd1 vccd1 _5481_/B sky130_fd_sc_hd__xnor2_1
X_7216_ _7233_/A _7233_/B vssd1 vssd1 vccd1 vccd1 _7216_/Y sky130_fd_sc_hd__nand2_1
X_4428_ _4431_/A vssd1 vssd1 vccd1 vccd1 _4428_/Y sky130_fd_sc_hd__inv_2
X_8196_ _8196_/A _8283_/A vssd1 vssd1 vccd1 vccd1 _8196_/X sky130_fd_sc_hd__or2_1
XFILLER_98_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4359_ _4363_/A vssd1 vssd1 vccd1 vccd1 _4359_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7147_ _7147_/A _7147_/B _7167_/A vssd1 vssd1 vccd1 vccd1 _7148_/B sky130_fd_sc_hd__nor3_1
XFILLER_59_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7078_ _7078_/A _7078_/B vssd1 vssd1 vccd1 vccd1 _7078_/Y sky130_fd_sc_hd__nor2_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8813__80 vssd1 vssd1 vccd1 vccd1 _8813__80/HI _8922_/A sky130_fd_sc_hd__conb_1
XFILLER_73_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6029_ _6030_/A _5747_/B _6095_/A vssd1 vssd1 vccd1 vccd1 _6096_/A sky130_fd_sc_hd__a21oi_1
XFILLER_73_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6380_ _8681_/Q vssd1 vssd1 vccd1 vccd1 _6426_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5400_ _5400_/A _8656_/Q vssd1 vssd1 vccd1 vccd1 _5401_/B sky130_fd_sc_hd__or2b_1
X_5331_ _5331_/A vssd1 vssd1 vccd1 vccd1 _8643_/D sky130_fd_sc_hd__clkbuf_1
X_8050_ _8110_/A _8110_/B vssd1 vssd1 vccd1 vccd1 _8082_/A sky130_fd_sc_hd__xor2_1
X_7001_ _7328_/A _7001_/B vssd1 vssd1 vccd1 vccd1 _7329_/B sky130_fd_sc_hd__nor2_1
X_5262_ _8665_/Q _5258_/X _5261_/X _4651_/X vssd1 vssd1 vccd1 vccd1 _8623_/D sky130_fd_sc_hd__o211a_1
XFILLER_87_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5193_ _5193_/A _5193_/B vssd1 vssd1 vccd1 vccd1 _5209_/B sky130_fd_sc_hd__or2_1
XFILLER_68_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8883_ _8883_/A _4396_/Y vssd1 vssd1 vccd1 vccd1 io_out[20] sky130_fd_sc_hd__ebufn_8
X_7903_ _8054_/A _8071_/A _7903_/C vssd1 vssd1 vccd1 vccd1 _7903_/X sky130_fd_sc_hd__and3_1
XFILLER_70_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7834_ _7834_/A _7835_/B vssd1 vssd1 vccd1 vccd1 _8052_/A sky130_fd_sc_hd__or2_1
XFILLER_24_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7765_ _8610_/Q _8571_/A vssd1 vssd1 vccd1 vccd1 _7771_/A sky130_fd_sc_hd__or2b_2
X_6716_ _7348_/B _6694_/B _6804_/A _7172_/B _7254_/B vssd1 vssd1 vccd1 vccd1 _6716_/X
+ sky130_fd_sc_hd__a32o_1
X_4977_ _4977_/A _5127_/A vssd1 vssd1 vccd1 vccd1 _5172_/B sky130_fd_sc_hd__or2_1
XFILLER_11_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7696_ _7711_/A _7703_/B vssd1 vssd1 vccd1 vccd1 _7728_/A sky130_fd_sc_hd__nand2_2
X_6647_ _6710_/A vssd1 vssd1 vccd1 vccd1 _6980_/A sky130_fd_sc_hd__buf_2
X_6578_ _6588_/A _6578_/B vssd1 vssd1 vccd1 vccd1 _6734_/A sky130_fd_sc_hd__xnor2_2
X_8317_ _8317_/A _8317_/B vssd1 vssd1 vccd1 vccd1 _8383_/A sky130_fd_sc_hd__xnor2_2
XFILLER_3_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5529_ _6070_/B _5541_/A vssd1 vssd1 vccd1 vccd1 _5530_/A sky130_fd_sc_hd__or2_1
XFILLER_59_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8248_ _8473_/S _8247_/X _8152_/B _8152_/A vssd1 vssd1 vccd1 vccd1 _8277_/B sky130_fd_sc_hd__a2bb2o_1
X_8179_ _8179_/A _8179_/B vssd1 vssd1 vccd1 vccd1 _8180_/B sky130_fd_sc_hd__nand2_1
XFILLER_59_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4900_ _4900_/A _4900_/B _5087_/B vssd1 vssd1 vccd1 vccd1 _5238_/C sky130_fd_sc_hd__and3_1
XFILLER_52_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5880_ _5978_/A _5880_/B vssd1 vssd1 vccd1 vccd1 _5905_/A sky130_fd_sc_hd__and2_1
X_4831_ _5244_/B _5230_/B vssd1 vssd1 vccd1 vccd1 _5044_/B sky130_fd_sc_hd__or2_1
XFILLER_33_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7550_ _7550_/A _7550_/B _7550_/C vssd1 vssd1 vccd1 vccd1 _7551_/A sky130_fd_sc_hd__and3_1
X_4762_ _4762_/A vssd1 vssd1 vccd1 vccd1 _8615_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4693_ _4694_/A _4711_/A vssd1 vssd1 vccd1 vccd1 _4700_/A sky130_fd_sc_hd__nand2_1
X_6501_ _6493_/X _6500_/Y _8558_/A vssd1 vssd1 vccd1 vccd1 _8697_/D sky130_fd_sc_hd__a21o_1
X_7481_ _7481_/A _7481_/B vssd1 vssd1 vccd1 vccd1 _7482_/B sky130_fd_sc_hd__nand2_1
X_6432_ _8684_/Q _8683_/Q _6432_/C vssd1 vssd1 vccd1 vccd1 _6437_/C sky130_fd_sc_hd__and3_1
X_8102_ _8102_/A _8102_/B vssd1 vssd1 vccd1 vccd1 _8506_/A sky130_fd_sc_hd__nor2_2
X_6363_ _6364_/A _6364_/B vssd1 vssd1 vccd1 vccd1 _6363_/Y sky130_fd_sc_hd__nand2_1
X_5314_ _8639_/Q _8638_/Q _5314_/C vssd1 vssd1 vccd1 vccd1 _5322_/C sky130_fd_sc_hd__and3_1
XFILLER_88_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6294_ _6294_/A _6294_/B vssd1 vssd1 vccd1 vccd1 _6336_/A sky130_fd_sc_hd__xnor2_4
X_5245_ _5245_/A _5245_/B _5245_/C _5245_/D vssd1 vssd1 vccd1 vccd1 _5245_/X sky130_fd_sc_hd__or4_1
X_8033_ _8114_/A _8114_/B vssd1 vssd1 vccd1 vccd1 _8042_/A sky130_fd_sc_hd__xnor2_1
XFILLER_102_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5176_ _5218_/D _5174_/X _5175_/X vssd1 vssd1 vccd1 vccd1 _5177_/C sky130_fd_sc_hd__o21a_1
XFILLER_56_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8935_ _8935_/A _4457_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[34] sky130_fd_sc_hd__ebufn_8
XFILLER_83_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_5_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_101_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8866_ _8866_/A _4374_/Y vssd1 vssd1 vccd1 vccd1 io_out[3] sky130_fd_sc_hd__ebufn_8
XFILLER_64_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7817_ _7817_/A _7817_/B vssd1 vssd1 vccd1 vccd1 _7818_/B sky130_fd_sc_hd__nor2_1
XFILLER_61_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7748_ _7748_/A _7748_/B vssd1 vssd1 vccd1 vccd1 _7748_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_20_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7679_ _8731_/Q _8607_/Q vssd1 vssd1 vccd1 vccd1 _7681_/A sky130_fd_sc_hd__and2b_1
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5030_ _5030_/A vssd1 vssd1 vccd1 vccd1 _5096_/A sky130_fd_sc_hd__clkbuf_2
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6981_ _6730_/A _6730_/B _6848_/A _6848_/B _7332_/A vssd1 vssd1 vccd1 vccd1 _7031_/S
+ sky130_fd_sc_hd__a221o_1
XFILLER_80_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5932_ _5924_/A _5924_/B _5925_/A _5923_/A vssd1 vssd1 vccd1 vccd1 _6013_/A sky130_fd_sc_hd__a31o_1
X_8720_ _8732_/CLK _8720_/D vssd1 vssd1 vccd1 vccd1 _8720_/Q sky130_fd_sc_hd__dfxtp_1
X_8651_ _8677_/CLK _8651_/D vssd1 vssd1 vccd1 vccd1 _8651_/Q sky130_fd_sc_hd__dfxtp_1
X_5863_ _5970_/B _5863_/B vssd1 vssd1 vccd1 vccd1 _5863_/Y sky130_fd_sc_hd__nor2_1
X_4814_ _4845_/A _4845_/B _4845_/C _4848_/C vssd1 vssd1 vccd1 vccd1 _4827_/A sky130_fd_sc_hd__or4_4
X_7602_ _7602_/A vssd1 vssd1 vccd1 vccd1 _8720_/D sky130_fd_sc_hd__clkbuf_1
X_5794_ _5889_/A _5794_/B vssd1 vssd1 vccd1 vccd1 _5795_/B sky130_fd_sc_hd__xnor2_1
X_8582_ _8672_/CLK _8582_/D vssd1 vssd1 vccd1 vccd1 _8582_/Q sky130_fd_sc_hd__dfxtp_1
X_7533_ _7533_/A _7533_/B vssd1 vssd1 vccd1 vccd1 _7535_/B sky130_fd_sc_hd__nand2_1
X_4745_ _5265_/A vssd1 vssd1 vccd1 vccd1 _5263_/B sky130_fd_sc_hd__clkbuf_2
X_7464_ _7390_/A _7390_/B _7463_/Y vssd1 vssd1 vccd1 vccd1 _7465_/B sky130_fd_sc_hd__o21a_1
X_4676_ _4942_/A vssd1 vssd1 vccd1 vccd1 _5143_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6415_ _6415_/A vssd1 vssd1 vccd1 vccd1 _8678_/D sky130_fd_sc_hd__clkbuf_1
X_7395_ _7395_/A _7395_/B vssd1 vssd1 vccd1 vccd1 _7395_/X sky130_fd_sc_hd__or2_1
X_6346_ _6346_/A _6353_/B vssd1 vssd1 vccd1 vccd1 _6347_/B sky130_fd_sc_hd__nand2_1
XFILLER_103_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6277_ _6278_/A _6278_/B vssd1 vssd1 vccd1 vccd1 _6277_/Y sky130_fd_sc_hd__nor2_1
X_8016_ _8019_/A _8015_/C _8015_/A vssd1 vssd1 vccd1 vccd1 _8017_/C sky130_fd_sc_hd__o21ai_1
XFILLER_102_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5228_ _5102_/B _5227_/X _5243_/A vssd1 vssd1 vccd1 vccd1 _5229_/D sky130_fd_sc_hd__o21a_1
XFILLER_29_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5159_ _5154_/A _5175_/C _5106_/C _5172_/B _5200_/C vssd1 vssd1 vccd1 vccd1 _5159_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_29_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8918_ _8918_/A _4436_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[17] sky130_fd_sc_hd__ebufn_8
X_8849_ _8849_/A _4355_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[18] sky130_fd_sc_hd__ebufn_8
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8774__41 vssd1 vssd1 vccd1 vccd1 _8774__41/HI _8869_/A sky130_fd_sc_hd__conb_1
XFILLER_28_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4530_ _4845_/A vssd1 vssd1 vccd1 vccd1 _4839_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_7_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4461_ _4461_/A vssd1 vssd1 vccd1 vccd1 _4461_/Y sky130_fd_sc_hd__inv_2
X_7180_ _7187_/A _7187_/B _7179_/X vssd1 vssd1 vccd1 vccd1 _7225_/A sky130_fd_sc_hd__a21oi_1
X_6200_ _6200_/A _6007_/B vssd1 vssd1 vccd1 vccd1 _6201_/B sky130_fd_sc_hd__or2b_1
X_4392_ _4394_/A vssd1 vssd1 vccd1 vccd1 _4392_/Y sky130_fd_sc_hd__inv_2
X_6131_ _6316_/B _5831_/X _6119_/B _6133_/B _6130_/A vssd1 vssd1 vccd1 vccd1 _6146_/B
+ sky130_fd_sc_hd__a41o_1
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6062_ _6157_/A _6303_/B vssd1 vssd1 vccd1 vccd1 _6062_/Y sky130_fd_sc_hd__xnor2_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5013_ _5016_/A _5155_/B vssd1 vssd1 vccd1 vccd1 _5022_/B sky130_fd_sc_hd__or2_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6964_ _6964_/A _6964_/B _6964_/C vssd1 vssd1 vccd1 vccd1 _6967_/A sky130_fd_sc_hd__nand3_1
XFILLER_53_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6895_ _7002_/A vssd1 vssd1 vccd1 vccd1 _7327_/A sky130_fd_sc_hd__clkbuf_2
X_8703_ _8703_/CLK _8703_/D vssd1 vssd1 vccd1 vccd1 _8703_/Q sky130_fd_sc_hd__dfxtp_1
X_5915_ _5936_/A _5936_/B vssd1 vssd1 vccd1 vccd1 _5916_/B sky130_fd_sc_hd__xor2_1
X_8634_ _8710_/CLK _8634_/D vssd1 vssd1 vccd1 vccd1 _8634_/Q sky130_fd_sc_hd__dfxtp_1
X_5846_ _5846_/A _5846_/B vssd1 vssd1 vccd1 vccd1 _5847_/B sky130_fd_sc_hd__nand2_1
XFILLER_61_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8565_ _8577_/S _8565_/B vssd1 vssd1 vccd1 vccd1 _8565_/X sky130_fd_sc_hd__and2_1
XFILLER_21_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5777_ _5788_/B _5777_/B vssd1 vssd1 vccd1 vccd1 _5802_/A sky130_fd_sc_hd__xnor2_1
X_7516_ _7516_/A _7516_/B vssd1 vssd1 vccd1 vccd1 _7517_/B sky130_fd_sc_hd__nand2_1
X_4728_ _4728_/A vssd1 vssd1 vccd1 vccd1 _8609_/D sky130_fd_sc_hd__clkbuf_1
X_8496_ _8496_/A _8496_/B _8496_/C vssd1 vssd1 vccd1 vccd1 _8496_/X sky130_fd_sc_hd__and3_1
X_7447_ _7455_/B _7447_/B _7447_/C _7447_/D vssd1 vssd1 vccd1 vccd1 _7449_/A sky130_fd_sc_hd__nand4_1
X_4659_ _4845_/C _8612_/Q _4898_/A vssd1 vssd1 vccd1 vccd1 _5047_/A sky130_fd_sc_hd__or3_4
XFILLER_101_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7378_ _7378_/A _7378_/B _7378_/C _7378_/D vssd1 vssd1 vccd1 vccd1 _7378_/Y sky130_fd_sc_hd__nor4_2
XFILLER_103_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6329_ _6336_/A _6336_/B _6331_/A _6329_/D vssd1 vssd1 vccd1 vccd1 _6329_/X sky130_fd_sc_hd__or4_1
XFILLER_76_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5700_ _5698_/X _5582_/B _5699_/Y vssd1 vssd1 vccd1 vccd1 _5721_/A sky130_fd_sc_hd__a21boi_2
X_6680_ _7254_/B _6957_/B _7169_/B _6655_/A vssd1 vssd1 vccd1 vccd1 _6702_/B sky130_fd_sc_hd__a22o_1
X_5631_ _5739_/B vssd1 vssd1 vccd1 vccd1 _5746_/B sky130_fd_sc_hd__clkbuf_2
X_8350_ _8350_/A _8359_/B vssd1 vssd1 vccd1 vccd1 _8351_/B sky130_fd_sc_hd__xnor2_1
X_5562_ _5998_/A _5992_/A vssd1 vssd1 vccd1 vccd1 _5571_/A sky130_fd_sc_hd__nor2_1
X_7301_ _7041_/A _7041_/B _7300_/X vssd1 vssd1 vccd1 vccd1 _7390_/A sky130_fd_sc_hd__a21oi_1
X_4513_ _8605_/Q vssd1 vssd1 vccd1 vccd1 _7695_/B sky130_fd_sc_hd__clkbuf_4
X_8281_ _8281_/A _8281_/B vssd1 vssd1 vccd1 vccd1 _8281_/Y sky130_fd_sc_hd__nor2_1
X_7232_ _7232_/A _7232_/B vssd1 vssd1 vccd1 vccd1 _7250_/A sky130_fd_sc_hd__xor2_1
X_5493_ _5493_/A _5493_/B _5493_/C vssd1 vssd1 vccd1 vccd1 _5506_/A sky130_fd_sc_hd__nand3_1
X_4444_ _4456_/A vssd1 vssd1 vccd1 vccd1 _4449_/A sky130_fd_sc_hd__clkbuf_2
X_4375_ _4375_/A vssd1 vssd1 vccd1 vccd1 _4375_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7163_ _7291_/A _7163_/B vssd1 vssd1 vccd1 vccd1 _7292_/B sky130_fd_sc_hd__xnor2_1
XFILLER_98_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7094_ _7105_/A _7105_/C _7105_/B vssd1 vssd1 vccd1 vccd1 _7097_/A sky130_fd_sc_hd__a21bo_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6114_ _6143_/A _6113_/C _6113_/A vssd1 vssd1 vccd1 vccd1 _6115_/B sky130_fd_sc_hd__a21o_1
XFILLER_100_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6045_ _6046_/A _6045_/B _6044_/X vssd1 vssd1 vccd1 vccd1 _6046_/B sky130_fd_sc_hd__nor3b_1
XFILLER_100_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7996_ _8063_/A vssd1 vssd1 vccd1 vccd1 _8072_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_26_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6947_ _7119_/B _7119_/A vssd1 vssd1 vccd1 vccd1 _6947_/X sky130_fd_sc_hd__or2b_1
XFILLER_54_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6878_ _7352_/A _7352_/C vssd1 vssd1 vccd1 vccd1 _6879_/A sky130_fd_sc_hd__nor2_1
XFILLER_34_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8617_ _8733_/CLK _8617_/D vssd1 vssd1 vccd1 vccd1 _8617_/Q sky130_fd_sc_hd__dfxtp_2
X_5829_ _5829_/A _5829_/B vssd1 vssd1 vccd1 vccd1 _5854_/B sky130_fd_sc_hd__xor2_1
X_8548_ _8548_/A _8548_/B vssd1 vssd1 vccd1 vccd1 _8550_/A sky130_fd_sc_hd__nor2_1
X_8479_ _8479_/A _8479_/B vssd1 vssd1 vccd1 vccd1 _8484_/A sky130_fd_sc_hd__xnor2_1
XFILLER_78_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8744__11 vssd1 vssd1 vccd1 vccd1 _8744__11/HI _8839_/A sky130_fd_sc_hd__conb_1
XFILLER_60_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7850_ _7850_/A _7850_/B vssd1 vssd1 vccd1 vccd1 _7940_/B sky130_fd_sc_hd__or2_1
XFILLER_36_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6801_ _6801_/A _6907_/B vssd1 vssd1 vccd1 vccd1 _6802_/B sky130_fd_sc_hd__xnor2_1
XFILLER_90_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4993_ _4993_/A vssd1 vssd1 vccd1 vccd1 _5227_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7781_ _7781_/A _7854_/C vssd1 vssd1 vccd1 vccd1 _7792_/A sky130_fd_sc_hd__xnor2_1
X_6732_ _7332_/B vssd1 vssd1 vccd1 vccd1 _7054_/B sky130_fd_sc_hd__clkbuf_2
X_6663_ _6663_/A _6663_/B vssd1 vssd1 vccd1 vccd1 _6677_/A sky130_fd_sc_hd__nand2_2
X_5614_ _5641_/A _5614_/B vssd1 vssd1 vccd1 vccd1 _5813_/A sky130_fd_sc_hd__xnor2_2
X_8402_ _8402_/A _8402_/B vssd1 vssd1 vccd1 vccd1 _8404_/C sky130_fd_sc_hd__xnor2_1
X_6594_ _8715_/Q vssd1 vssd1 vccd1 vccd1 _7548_/A sky130_fd_sc_hd__clkinv_2
X_5545_ _6020_/A _5993_/A _5713_/A vssd1 vssd1 vccd1 vccd1 _5545_/Y sky130_fd_sc_hd__a21oi_1
X_8333_ _8396_/A _8396_/B vssd1 vssd1 vccd1 vccd1 _8397_/B sky130_fd_sc_hd__xor2_1
X_8264_ _8499_/A _8499_/B vssd1 vssd1 vccd1 vccd1 _8264_/Y sky130_fd_sc_hd__xnor2_1
X_5476_ _5517_/A vssd1 vssd1 vccd1 vccd1 _5566_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7215_ _7215_/A _7215_/B vssd1 vssd1 vccd1 vccd1 _7233_/B sky130_fd_sc_hd__xnor2_1
X_4427_ _4431_/A vssd1 vssd1 vccd1 vccd1 _4427_/Y sky130_fd_sc_hd__inv_2
X_8195_ _8195_/A _8195_/B vssd1 vssd1 vccd1 vccd1 _8199_/A sky130_fd_sc_hd__and2_1
X_7146_ _7146_/A _7146_/B vssd1 vssd1 vccd1 vccd1 _7177_/A sky130_fd_sc_hd__xor2_1
X_4358_ _4370_/A vssd1 vssd1 vccd1 vccd1 _4363_/A sky130_fd_sc_hd__clkbuf_2
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7077_ _7078_/A _7078_/B vssd1 vssd1 vccd1 vccd1 _7138_/B sky130_fd_sc_hd__xor2_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6028_ _6028_/A _6028_/B vssd1 vssd1 vccd1 vccd1 _6095_/A sky130_fd_sc_hd__nor2_1
XFILLER_104_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7979_ _8024_/B _7978_/C _7978_/A vssd1 vssd1 vccd1 vccd1 _7980_/C sky130_fd_sc_hd__a21o_1
XFILLER_42_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5330_ _5332_/B _5330_/B _5362_/A vssd1 vssd1 vccd1 vccd1 _5331_/A sky130_fd_sc_hd__and3b_1
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5261_ _8623_/Q _5263_/B vssd1 vssd1 vccd1 vccd1 _5261_/X sky130_fd_sc_hd__or2_1
Xclkbuf_4_7_0_wb_clk_i clkbuf_4_7_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _8734_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_102_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7000_ _7000_/A _7000_/B vssd1 vssd1 vccd1 vccd1 _7001_/B sky130_fd_sc_hd__and2_1
X_5192_ _5192_/A _5192_/B _5200_/B _5192_/D vssd1 vssd1 vccd1 vccd1 _5192_/X sky130_fd_sc_hd__or4_1
XFILLER_83_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7902_ _8065_/B vssd1 vssd1 vccd1 vccd1 _8071_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_70_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8882_ _8882_/A _4394_/Y vssd1 vssd1 vccd1 vccd1 io_out[19] sky130_fd_sc_hd__ebufn_8
XFILLER_36_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7833_ _7833_/A _7833_/B vssd1 vssd1 vccd1 vccd1 _7847_/A sky130_fd_sc_hd__xnor2_1
X_7764_ _8124_/A _7857_/C vssd1 vssd1 vccd1 vccd1 _7780_/A sky130_fd_sc_hd__xnor2_1
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4976_ _5164_/C vssd1 vssd1 vccd1 vccd1 _5009_/B sky130_fd_sc_hd__clkbuf_2
X_6715_ _6715_/A vssd1 vssd1 vccd1 vccd1 _7348_/B sky130_fd_sc_hd__clkbuf_2
X_7695_ _7695_/A _7695_/B vssd1 vssd1 vccd1 vccd1 _7703_/B sky130_fd_sc_hd__nand2_1
X_6646_ _6589_/A _7000_/A _6872_/A vssd1 vssd1 vccd1 vccd1 _6710_/A sky130_fd_sc_hd__mux2_1
X_6577_ _7128_/A _6711_/A vssd1 vssd1 vccd1 vccd1 _7275_/A sky130_fd_sc_hd__or2_2
X_8316_ _8316_/A _8316_/B vssd1 vssd1 vccd1 vccd1 _8317_/B sky130_fd_sc_hd__xor2_1
X_5528_ _5493_/A _5491_/B _5493_/C _5489_/X vssd1 vssd1 vccd1 vccd1 _5541_/A sky130_fd_sc_hd__a31o_1
XFILLER_3_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8247_ _8308_/A _8247_/B vssd1 vssd1 vccd1 vccd1 _8247_/X sky130_fd_sc_hd__or2_1
X_5459_ _5475_/A _5475_/B vssd1 vssd1 vccd1 vccd1 _5780_/A sky130_fd_sc_hd__xor2_2
X_8178_ _8178_/A _8178_/B vssd1 vssd1 vccd1 vccd1 _8179_/B sky130_fd_sc_hd__or2_1
XFILLER_86_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7129_ _7133_/A _7132_/A vssd1 vssd1 vccd1 vccd1 _7131_/A sky130_fd_sc_hd__nand2_1
XFILLER_86_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4830_ _4830_/A _4849_/B vssd1 vssd1 vccd1 vccd1 _5230_/B sky130_fd_sc_hd__nor2_2
XFILLER_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4761_ _8544_/A _4761_/B vssd1 vssd1 vccd1 vccd1 _4762_/A sky130_fd_sc_hd__and2_1
X_6500_ _6500_/A _6500_/B vssd1 vssd1 vccd1 vccd1 _6500_/Y sky130_fd_sc_hd__nand2_1
X_4692_ _4692_/A vssd1 vssd1 vccd1 vccd1 _4694_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7480_ _7480_/A _7480_/B vssd1 vssd1 vccd1 vccd1 _7480_/X sky130_fd_sc_hd__xor2_1
X_6431_ _6431_/A _6431_/B vssd1 vssd1 vccd1 vccd1 _8683_/D sky130_fd_sc_hd__nor2_1
X_6362_ _6355_/B _6356_/A _6354_/B _6355_/A vssd1 vssd1 vccd1 vccd1 _6364_/B sky130_fd_sc_hd__o211a_1
X_5313_ _6466_/B _5314_/C _5312_/Y vssd1 vssd1 vccd1 vccd1 _8638_/D sky130_fd_sc_hd__a21oi_1
X_8101_ _8101_/A _8102_/B _8503_/A _8100_/X vssd1 vssd1 vccd1 vccd1 _8506_/B sky130_fd_sc_hd__or4bb_2
X_6293_ _6293_/A _6293_/B vssd1 vssd1 vccd1 vccd1 _6294_/B sky130_fd_sc_hd__xnor2_4
XFILLER_88_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5244_ _5244_/A _5244_/B _5244_/C vssd1 vssd1 vccd1 vccd1 _5244_/X sky130_fd_sc_hd__or3_1
X_8032_ _8044_/A _8032_/B vssd1 vssd1 vccd1 vccd1 _8114_/B sky130_fd_sc_hd__xnor2_1
X_5175_ _5175_/A _5175_/B _5175_/C _5175_/D vssd1 vssd1 vccd1 vccd1 _5175_/X sky130_fd_sc_hd__or4_1
XFILLER_56_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8934_ _8934_/A _4455_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[33] sky130_fd_sc_hd__ebufn_8
X_8865_ _8865_/A _4373_/Y vssd1 vssd1 vccd1 vccd1 io_out[2] sky130_fd_sc_hd__ebufn_8
XFILLER_71_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7816_ _7815_/B _7901_/A vssd1 vssd1 vccd1 vccd1 _7817_/B sky130_fd_sc_hd__and2b_1
XFILLER_101_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4959_ _5153_/A _5111_/A _5136_/B _5244_/C _4914_/X vssd1 vssd1 vccd1 vccd1 _4959_/X
+ sky130_fd_sc_hd__o32a_1
X_7747_ _8063_/A _7798_/B _7813_/B _7746_/X vssd1 vssd1 vccd1 vccd1 _7748_/B sky130_fd_sc_hd__a31oi_2
X_7678_ _7769_/A _7678_/B vssd1 vssd1 vccd1 vccd1 _7759_/A sky130_fd_sc_hd__nor2_4
X_6629_ _8700_/Q _5591_/A vssd1 vssd1 vccd1 vccd1 _6631_/A sky130_fd_sc_hd__or2b_1
XFILLER_20_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6980_ _6980_/A _7336_/S vssd1 vssd1 vccd1 vccd1 _6984_/A sky130_fd_sc_hd__nor2_1
XFILLER_93_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5931_ _5928_/A _5928_/B _5930_/Y vssd1 vssd1 vccd1 vccd1 _6160_/A sky130_fd_sc_hd__a21oi_1
XFILLER_25_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8650_ _8677_/CLK _8650_/D vssd1 vssd1 vccd1 vccd1 _8650_/Q sky130_fd_sc_hd__dfxtp_1
X_5862_ _5970_/B _5863_/B vssd1 vssd1 vccd1 vccd1 _5862_/Y sky130_fd_sc_hd__nand2_1
XFILLER_33_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4813_ _4879_/A vssd1 vssd1 vccd1 vccd1 _4919_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_21_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7601_ _8544_/A _7601_/B vssd1 vssd1 vccd1 vccd1 _7602_/A sky130_fd_sc_hd__and2_1
X_5793_ _5998_/A _5884_/B vssd1 vssd1 vccd1 vccd1 _5889_/A sky130_fd_sc_hd__or2_1
X_8581_ _8672_/CLK _8581_/D vssd1 vssd1 vccd1 vccd1 _8581_/Q sky130_fd_sc_hd__dfxtp_1
X_7532_ _7546_/A _7532_/B vssd1 vssd1 vccd1 vccd1 _7533_/B sky130_fd_sc_hd__or2_1
X_4744_ _4763_/A _4752_/A vssd1 vssd1 vccd1 vccd1 _5265_/A sky130_fd_sc_hd__and2_1
X_7463_ _7463_/A _7463_/B vssd1 vssd1 vccd1 vccd1 _7463_/Y sky130_fd_sc_hd__nand2_1
X_4675_ _5244_/A vssd1 vssd1 vccd1 vccd1 _4942_/A sky130_fd_sc_hd__buf_2
X_6414_ _6418_/C _6414_/B _6457_/B vssd1 vssd1 vccd1 vccd1 _6415_/A sky130_fd_sc_hd__and3b_1
X_7394_ _7397_/A _7397_/B vssd1 vssd1 vccd1 vccd1 _7394_/X sky130_fd_sc_hd__xor2_1
X_6345_ _6346_/A _6353_/B vssd1 vssd1 vccd1 vccd1 _6355_/A sky130_fd_sc_hd__or2_1
X_6276_ _6276_/A _6276_/B vssd1 vssd1 vccd1 vccd1 _6280_/A sky130_fd_sc_hd__xnor2_1
XFILLER_88_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5227_ _5227_/A _5227_/B _5227_/C _5227_/D vssd1 vssd1 vccd1 vccd1 _5227_/X sky130_fd_sc_hd__or4_1
X_8015_ _8015_/A _8019_/A _8015_/C vssd1 vssd1 vccd1 vccd1 _8017_/B sky130_fd_sc_hd__or3_1
XFILLER_88_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5158_ _4707_/A _5152_/X _5157_/X _5096_/A _5080_/Y vssd1 vssd1 vccd1 vccd1 _5158_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_56_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5089_ _5130_/A _5091_/C _5238_/B _5089_/D vssd1 vssd1 vccd1 vccd1 _5089_/X sky130_fd_sc_hd__or4_1
XFILLER_56_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8917_ _8917_/A _4435_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[16] sky130_fd_sc_hd__ebufn_8
XFILLER_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8848_ _8848_/A _4354_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[17] sky130_fd_sc_hd__ebufn_8
XFILLER_72_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4460_ _4461_/A vssd1 vssd1 vccd1 vccd1 _4460_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4391_ _4394_/A vssd1 vssd1 vccd1 vccd1 _4391_/Y sky130_fd_sc_hd__inv_2
X_6130_ _6130_/A _6130_/B vssd1 vssd1 vccd1 vccd1 _6133_/B sky130_fd_sc_hd__nor2_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6061_ _6061_/A _6061_/B vssd1 vssd1 vccd1 vccd1 _6303_/B sky130_fd_sc_hd__nor2_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5012_ _5227_/A _5154_/B vssd1 vssd1 vccd1 vccd1 _5155_/B sky130_fd_sc_hd__or2_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6963_ _7361_/A _6962_/C _7355_/A vssd1 vssd1 vccd1 vccd1 _6964_/C sky130_fd_sc_hd__o21ai_1
XFILLER_81_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6894_ _6775_/A _6798_/Y _6722_/X _6893_/X vssd1 vssd1 vccd1 vccd1 _7002_/A sky130_fd_sc_hd__a211o_1
XFILLER_81_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8702_ _8703_/CLK _8702_/D vssd1 vssd1 vccd1 vccd1 _8702_/Q sky130_fd_sc_hd__dfxtp_1
X_5914_ _5746_/B _5970_/A _5816_/B _5819_/A _5819_/B vssd1 vssd1 vccd1 vccd1 _5936_/B
+ sky130_fd_sc_hd__a32o_1
X_8633_ _8734_/CLK _8633_/D vssd1 vssd1 vccd1 vccd1 _8633_/Q sky130_fd_sc_hd__dfxtp_1
X_5845_ _5845_/A _5845_/B vssd1 vssd1 vccd1 vccd1 _5846_/B sky130_fd_sc_hd__or2_1
XFILLER_22_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8564_ _8563_/A _8563_/C _8563_/B vssd1 vssd1 vccd1 vccd1 _8565_/B sky130_fd_sc_hd__o21ai_1
X_5776_ _5720_/A _5720_/B _5775_/Y vssd1 vssd1 vccd1 vccd1 _5801_/A sky130_fd_sc_hd__o21a_1
XFILLER_21_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7515_ _7516_/A _7516_/B vssd1 vssd1 vccd1 vccd1 _7515_/Y sky130_fd_sc_hd__nor2_1
X_4727_ _4727_/A _4727_/B _4730_/B vssd1 vssd1 vccd1 vccd1 _4728_/A sky130_fd_sc_hd__and3_1
XFILLER_21_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8495_ _8496_/B _8496_/C _8496_/A vssd1 vssd1 vccd1 vccd1 _8495_/Y sky130_fd_sc_hd__a21oi_1
X_7446_ _6880_/X _6958_/B _7352_/X _7454_/B vssd1 vssd1 vccd1 vccd1 _7450_/A sky130_fd_sc_hd__o211ai_2
X_4658_ _4845_/A _4845_/B vssd1 vssd1 vccd1 vccd1 _4898_/A sky130_fd_sc_hd__nand2_2
X_7377_ _7376_/A _7376_/B _7376_/C vssd1 vssd1 vccd1 vccd1 _7378_/D sky130_fd_sc_hd__a21oi_1
XFILLER_89_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4589_ _8582_/Q _8581_/Q _8583_/Q vssd1 vssd1 vccd1 vccd1 _4598_/C sky130_fd_sc_hd__and3_1
X_6328_ _6332_/B _6332_/C vssd1 vssd1 vccd1 vccd1 _6329_/D sky130_fd_sc_hd__and2_1
XFILLER_67_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6259_ _6259_/A _6259_/B vssd1 vssd1 vccd1 vccd1 _6260_/B sky130_fd_sc_hd__xnor2_1
XFILLER_103_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5630_ _5630_/A _5630_/B vssd1 vssd1 vccd1 vccd1 _5739_/B sky130_fd_sc_hd__xnor2_2
X_5561_ _5709_/A vssd1 vssd1 vccd1 vccd1 _5893_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_31_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4512_ _4512_/A vssd1 vssd1 vccd1 vccd1 _8875_/A sky130_fd_sc_hd__buf_2
X_7300_ _7040_/B _7300_/B vssd1 vssd1 vccd1 vccd1 _7300_/X sky130_fd_sc_hd__and2b_1
X_8280_ _8515_/B _8243_/B _8246_/B _8279_/Y vssd1 vssd1 vccd1 vccd1 _8375_/B sky130_fd_sc_hd__a31o_1
X_5492_ _5470_/A _6598_/A _5475_/A _5475_/B _5447_/A vssd1 vssd1 vccd1 vccd1 _5493_/C
+ sky130_fd_sc_hd__a221o_1
X_7231_ _7231_/A vssd1 vssd1 vccd1 vccd1 _7479_/B sky130_fd_sc_hd__inv_2
XFILLER_7_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4443_ _4443_/A vssd1 vssd1 vccd1 vccd1 _4443_/Y sky130_fd_sc_hd__inv_2
X_4374_ _4375_/A vssd1 vssd1 vccd1 vccd1 _4374_/Y sky130_fd_sc_hd__inv_2
X_7162_ _7162_/A _7162_/B vssd1 vssd1 vccd1 vccd1 _7163_/B sky130_fd_sc_hd__xor2_1
X_7093_ _7101_/A _7101_/B _7093_/C vssd1 vssd1 vccd1 vccd1 _7105_/B sky130_fd_sc_hd__nand3_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6113_ _6113_/A _6143_/A _6113_/C vssd1 vssd1 vccd1 vccd1 _6143_/B sky130_fd_sc_hd__nand3_1
XFILLER_98_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6044_ _6051_/A _6044_/B vssd1 vssd1 vccd1 vccd1 _6044_/X sky130_fd_sc_hd__and2_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7995_ _8078_/A _8078_/B vssd1 vssd1 vccd1 vccd1 _8079_/A sky130_fd_sc_hd__xnor2_1
X_6946_ _6863_/A _6863_/B _6945_/X vssd1 vssd1 vccd1 vccd1 _7119_/A sky130_fd_sc_hd__a21bo_1
XFILLER_54_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6877_ _6890_/A vssd1 vssd1 vccd1 vccd1 _7352_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_8616_ _8733_/CLK _8616_/D vssd1 vssd1 vccd1 vccd1 _8616_/Q sky130_fd_sc_hd__dfxtp_4
X_5828_ _5922_/B _5828_/B vssd1 vssd1 vccd1 vccd1 _5829_/B sky130_fd_sc_hd__nor2_1
XFILLER_22_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5759_ _5941_/B _6273_/S _5962_/A vssd1 vssd1 vccd1 vccd1 _5763_/A sky130_fd_sc_hd__o21ai_1
X_8547_ _8547_/A _8560_/B vssd1 vssd1 vccd1 vccd1 _8548_/B sky130_fd_sc_hd__and2_1
X_8478_ _8478_/A _8478_/B vssd1 vssd1 vccd1 vccd1 _8479_/B sky130_fd_sc_hd__xnor2_1
X_7429_ _7429_/A _7429_/B vssd1 vssd1 vccd1 vccd1 _7461_/A sky130_fd_sc_hd__nor2_1
XFILLER_1_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6800_ _6800_/A _6999_/A vssd1 vssd1 vccd1 vccd1 _6907_/B sky130_fd_sc_hd__xor2_1
XFILLER_84_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4992_ _5207_/A _5245_/D _5164_/D vssd1 vssd1 vccd1 vccd1 _4992_/X sky130_fd_sc_hd__or3_1
X_7780_ _7780_/A _7780_/B vssd1 vssd1 vccd1 vccd1 _7854_/C sky130_fd_sc_hd__xor2_1
XFILLER_23_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6731_ _6829_/A vssd1 vssd1 vccd1 vccd1 _7332_/B sky130_fd_sc_hd__clkbuf_2
X_6662_ _6670_/B vssd1 vssd1 vccd1 vccd1 _6972_/C sky130_fd_sc_hd__buf_2
X_8401_ _8401_/A _8401_/B vssd1 vssd1 vccd1 vccd1 _8402_/B sky130_fd_sc_hd__xor2_1
X_5613_ _5610_/X _5619_/A _5619_/B _5621_/B vssd1 vssd1 vccd1 vccd1 _5614_/B sky130_fd_sc_hd__a31o_2
X_6593_ _6593_/A _6593_/B vssd1 vssd1 vccd1 vccd1 _7280_/A sky130_fd_sc_hd__nand2_4
X_8332_ _8410_/B _8332_/B vssd1 vssd1 vccd1 vccd1 _8396_/B sky130_fd_sc_hd__xor2_1
X_5544_ _6070_/B _5992_/B vssd1 vssd1 vccd1 vccd1 _5713_/A sky130_fd_sc_hd__nor2_1
X_8263_ _8430_/A _8430_/B vssd1 vssd1 vccd1 vccd1 _8499_/B sky130_fd_sc_hd__xor2_2
X_5475_ _5475_/A _5475_/B vssd1 vssd1 vccd1 vccd1 _5517_/A sky130_fd_sc_hd__xnor2_1
X_7214_ _7220_/A _7220_/B vssd1 vssd1 vccd1 vccd1 _7215_/B sky130_fd_sc_hd__xor2_1
X_4426_ _4432_/A vssd1 vssd1 vccd1 vccd1 _4431_/A sky130_fd_sc_hd__buf_6
X_8194_ _8402_/A vssd1 vssd1 vccd1 vccd1 _8195_/A sky130_fd_sc_hd__inv_2
X_7145_ _7145_/A _7145_/B vssd1 vssd1 vccd1 vccd1 _7146_/B sky130_fd_sc_hd__xnor2_2
XFILLER_98_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4357_ _4357_/A vssd1 vssd1 vccd1 vccd1 _4357_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7076_ _7102_/B _7076_/B vssd1 vssd1 vccd1 vccd1 _7078_/B sky130_fd_sc_hd__xor2_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6027_ _6038_/A _6035_/B vssd1 vssd1 vccd1 vccd1 _6027_/X sky130_fd_sc_hd__and2_1
XFILLER_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7978_ _7978_/A _8024_/B _7978_/C vssd1 vssd1 vccd1 vccd1 _8023_/A sky130_fd_sc_hd__nand3_1
XFILLER_54_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6929_ _7332_/B _6929_/B vssd1 vssd1 vccd1 vccd1 _6929_/Y sky130_fd_sc_hd__nor2_1
XFILLER_80_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_49_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8804__71 vssd1 vssd1 vccd1 vccd1 _8804__71/HI _8913_/A sky130_fd_sc_hd__conb_1
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5260_ _8664_/Q _5258_/X _5259_/X _4651_/X vssd1 vssd1 vccd1 vccd1 _8622_/D sky130_fd_sc_hd__o211a_1
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5191_ _5168_/X _5178_/X _5190_/X _4711_/B vssd1 vssd1 vccd1 vccd1 _5191_/X sky130_fd_sc_hd__a31o_1
XFILLER_95_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7901_ _7901_/A _7901_/B vssd1 vssd1 vccd1 vccd1 _8000_/A sky130_fd_sc_hd__nor2_1
X_8881_ _8881_/A _4393_/Y vssd1 vssd1 vccd1 vccd1 io_out[18] sky130_fd_sc_hd__ebufn_8
XFILLER_48_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7832_ _8101_/A _7832_/B vssd1 vssd1 vccd1 vccd1 _8533_/A sky130_fd_sc_hd__nand2_1
X_4975_ _5130_/A _5194_/A vssd1 vssd1 vccd1 vccd1 _5164_/C sky130_fd_sc_hd__nand2_2
X_7763_ _7779_/A _7763_/B vssd1 vssd1 vccd1 vccd1 _7857_/C sky130_fd_sc_hd__xnor2_1
X_6714_ _6768_/A _6768_/B vssd1 vssd1 vccd1 vccd1 _6769_/A sky130_fd_sc_hd__xnor2_1
X_7694_ _8729_/Q vssd1 vssd1 vccd1 vccd1 _7695_/A sky130_fd_sc_hd__inv_2
X_6645_ _6656_/B _6688_/A _6689_/A _6690_/A _6734_/A vssd1 vssd1 vccd1 vccd1 _6872_/A
+ sky130_fd_sc_hd__a311o_1
X_6576_ _6893_/C vssd1 vssd1 vccd1 vccd1 _6711_/A sky130_fd_sc_hd__clkbuf_2
X_8315_ _8460_/A _8386_/B vssd1 vssd1 vccd1 vccd1 _8316_/B sky130_fd_sc_hd__xnor2_1
X_5527_ _5540_/A _5527_/B vssd1 vssd1 vccd1 vccd1 _6070_/B sky130_fd_sc_hd__and2_2
X_8246_ _8483_/A _8246_/B vssd1 vssd1 vccd1 vccd1 _8277_/A sky130_fd_sc_hd__xnor2_1
X_5458_ _5480_/A _5480_/B _5477_/B _5457_/X _5455_/A vssd1 vssd1 vccd1 vccd1 _5475_/B
+ sky130_fd_sc_hd__a311o_4
X_4409_ _4413_/A vssd1 vssd1 vccd1 vccd1 _4409_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8177_ _8178_/A _8178_/B vssd1 vssd1 vccd1 vccd1 _8179_/A sky130_fd_sc_hd__nand2_1
X_5389_ _5389_/A _5389_/B vssd1 vssd1 vccd1 vccd1 _5389_/Y sky130_fd_sc_hd__nand2_1
X_7128_ _7128_/A _7128_/B vssd1 vssd1 vccd1 vccd1 _7132_/A sky130_fd_sc_hd__nor2_1
X_7059_ _7280_/A _7432_/A _7432_/B vssd1 vssd1 vccd1 vccd1 _7059_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_39_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4760_ _4758_/A _5285_/B _4844_/A _4759_/X vssd1 vssd1 vccd1 vccd1 _4761_/B sky130_fd_sc_hd__a22o_1
XFILLER_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4691_ _5205_/A vssd1 vssd1 vccd1 vccd1 _4692_/A sky130_fd_sc_hd__clkbuf_2
X_6430_ _8683_/Q _6432_/C _6423_/X vssd1 vssd1 vccd1 vccd1 _6431_/B sky130_fd_sc_hd__o21ai_1
X_6361_ _6366_/A _6361_/B vssd1 vssd1 vccd1 vccd1 _6364_/A sky130_fd_sc_hd__nand2_1
X_5312_ _6466_/B _5314_/C _5311_/X vssd1 vssd1 vccd1 vccd1 _5312_/Y sky130_fd_sc_hd__o21ai_1
X_8100_ _8017_/B _8017_/C _8017_/A vssd1 vssd1 vccd1 vccd1 _8100_/X sky130_fd_sc_hd__a21o_1
X_6292_ _6232_/A _6232_/B _6234_/B _6234_/A _6291_/Y vssd1 vssd1 vccd1 vccd1 _6293_/B
+ sky130_fd_sc_hd__a221oi_4
X_5243_ _5243_/A _5243_/B vssd1 vssd1 vccd1 vccd1 _5243_/X sky130_fd_sc_hd__and2_1
X_8031_ _8031_/A _8116_/A vssd1 vssd1 vccd1 vccd1 _8032_/B sky130_fd_sc_hd__xnor2_1
XFILLER_102_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5174_ _5237_/A _5171_/B _5175_/C _5173_/Y _5214_/A vssd1 vssd1 vccd1 vccd1 _5174_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_83_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8933_ _8933_/A _4454_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[32] sky130_fd_sc_hd__ebufn_8
XFILLER_83_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8864_ _8864_/A _4372_/Y vssd1 vssd1 vccd1 vccd1 io_out[1] sky130_fd_sc_hd__ebufn_8
X_8795__62 vssd1 vssd1 vccd1 vccd1 _8795__62/HI _8904_/A sky130_fd_sc_hd__conb_1
XFILLER_52_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7815_ _7901_/A _7815_/B vssd1 vssd1 vccd1 vccd1 _7817_/A sky130_fd_sc_hd__and2b_1
XFILLER_36_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4958_ _5091_/C _4958_/B vssd1 vssd1 vccd1 vccd1 _5244_/C sky130_fd_sc_hd__or2_2
X_7746_ _7835_/A _7813_/A _7835_/B _8145_/A vssd1 vssd1 vccd1 vccd1 _7746_/X sky130_fd_sc_hd__o22a_1
X_4889_ _4903_/B vssd1 vssd1 vccd1 vccd1 _4990_/A sky130_fd_sc_hd__clkbuf_2
X_7677_ _8733_/Q _7677_/B vssd1 vssd1 vccd1 vccd1 _7678_/B sky130_fd_sc_hd__and2_1
X_6628_ _7643_/B _8701_/Q vssd1 vssd1 vccd1 vccd1 _6659_/A sky130_fd_sc_hd__or2b_1
XFILLER_20_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6559_ _6559_/A _6559_/B vssd1 vssd1 vccd1 vccd1 _6835_/A sky130_fd_sc_hd__xnor2_4
XFILLER_3_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8229_ _8229_/A _8229_/B vssd1 vssd1 vccd1 vccd1 _8415_/B sky130_fd_sc_hd__nor2_2
XFILLER_59_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5930_ _5930_/A _5930_/B vssd1 vssd1 vccd1 vccd1 _5930_/Y sky130_fd_sc_hd__nor2_1
XFILLER_80_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5861_ _5861_/A _6196_/A vssd1 vssd1 vccd1 vccd1 _5869_/A sky130_fd_sc_hd__nand2_1
X_7600_ _7599_/Y _7596_/B _8543_/S vssd1 vssd1 vccd1 vccd1 _7601_/B sky130_fd_sc_hd__mux2_1
X_4812_ _4885_/B _4830_/A vssd1 vssd1 vccd1 vccd1 _4979_/A sky130_fd_sc_hd__nor2_2
XFILLER_61_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5792_ _5872_/A _5792_/B vssd1 vssd1 vccd1 vccd1 _5796_/A sky130_fd_sc_hd__nand2_1
X_8580_ _7876_/A _8578_/Y _8579_/Y vssd1 vssd1 vccd1 vccd1 _8735_/D sky130_fd_sc_hd__a21oi_1
X_7531_ _7546_/A _7532_/B vssd1 vssd1 vccd1 vccd1 _7533_/A sky130_fd_sc_hd__nand2_1
X_4743_ _4848_/B _4834_/C vssd1 vssd1 vccd1 vccd1 _4828_/C sky130_fd_sc_hd__nand2_1
XFILLER_21_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7462_ _7462_/A _7462_/B vssd1 vssd1 vccd1 vccd1 _7466_/A sky130_fd_sc_hd__xnor2_2
X_6413_ _8678_/Q _6413_/B vssd1 vssd1 vccd1 vccd1 _6414_/B sky130_fd_sc_hd__or2_1
X_4674_ _8603_/Q vssd1 vssd1 vccd1 vccd1 _5244_/A sky130_fd_sc_hd__inv_2
X_7393_ _7392_/A _7052_/B _7050_/Y vssd1 vssd1 vccd1 vccd1 _7397_/B sky130_fd_sc_hd__a21o_1
X_6344_ _6341_/A _5397_/X _5398_/X _6343_/Y vssd1 vssd1 vccd1 vccd1 _8669_/D sky130_fd_sc_hd__a22o_1
XFILLER_103_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6275_ _6275_/A _6275_/B vssd1 vssd1 vccd1 vccd1 _6276_/B sky130_fd_sc_hd__xnor2_1
XFILLER_102_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5226_ _5226_/A _5226_/B _5227_/B _5226_/D vssd1 vssd1 vccd1 vccd1 _5226_/X sky130_fd_sc_hd__or4_1
X_8014_ _8021_/B _8012_/X _7936_/A _7938_/A vssd1 vssd1 vccd1 vccd1 _8015_/C sky130_fd_sc_hd__a211oi_1
XFILLER_102_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5157_ _4702_/A _5015_/X _5153_/X _5156_/X _4694_/A vssd1 vssd1 vccd1 vccd1 _5157_/X
+ sky130_fd_sc_hd__o311a_1
X_5088_ _5200_/B _5119_/A _5199_/A vssd1 vssd1 vccd1 vccd1 _5089_/D sky130_fd_sc_hd__o21a_1
X_8916_ _8916_/A _4434_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[15] sky130_fd_sc_hd__ebufn_8
XFILLER_72_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8847_ _8847_/A _4353_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[16] sky130_fd_sc_hd__ebufn_8
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7729_ _7773_/A vssd1 vssd1 vccd1 vccd1 _8321_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_4_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4390_ _4394_/A vssd1 vssd1 vccd1 vccd1 _4390_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6060_ _6060_/A _6060_/B _6060_/C vssd1 vssd1 vccd1 vccd1 _6061_/B sky130_fd_sc_hd__nor3_1
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5011_ _5084_/C vssd1 vssd1 vccd1 vccd1 _5229_/B sky130_fd_sc_hd__clkbuf_2
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6962_ _7371_/A _7361_/A _6962_/C vssd1 vssd1 vccd1 vccd1 _6964_/B sky130_fd_sc_hd__or3_1
XFILLER_81_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8765__32 vssd1 vssd1 vccd1 vccd1 _8765__32/HI _8860_/A sky130_fd_sc_hd__conb_1
X_6893_ _6773_/X _6893_/B _6893_/C vssd1 vssd1 vccd1 vccd1 _6893_/X sky130_fd_sc_hd__and3b_1
X_8701_ _8733_/CLK _8701_/D vssd1 vssd1 vccd1 vccd1 _8701_/Q sky130_fd_sc_hd__dfxtp_1
X_5913_ _6242_/A _5913_/B vssd1 vssd1 vccd1 vccd1 _5936_/A sky130_fd_sc_hd__xnor2_1
X_8632_ _8734_/CLK _8632_/D vssd1 vssd1 vccd1 vccd1 _8632_/Q sky130_fd_sc_hd__dfxtp_1
X_5844_ _5845_/A _5845_/B vssd1 vssd1 vccd1 vccd1 _5846_/A sky130_fd_sc_hd__nand2_1
XFILLER_22_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8563_ _8563_/A _8563_/B _8563_/C vssd1 vssd1 vccd1 vccd1 _8577_/S sky130_fd_sc_hd__or3_1
X_7514_ _7514_/A _8696_/Q vssd1 vssd1 vccd1 vccd1 _7516_/B sky130_fd_sc_hd__xor2_1
X_5775_ _5775_/A _5775_/B vssd1 vssd1 vccd1 vccd1 _5775_/Y sky130_fd_sc_hd__nand2_1
X_4726_ _4801_/B _4726_/B vssd1 vssd1 vccd1 vccd1 _4730_/B sky130_fd_sc_hd__nand2_1
X_8494_ _8493_/A _8493_/B _8493_/C vssd1 vssd1 vccd1 vccd1 _8512_/B sky130_fd_sc_hd__a21oi_1
X_7445_ _7445_/A _7445_/B vssd1 vssd1 vccd1 vccd1 _7451_/A sky130_fd_sc_hd__xnor2_1
X_4657_ _5153_/A vssd1 vssd1 vccd1 vccd1 _4661_/A sky130_fd_sc_hd__clkbuf_2
X_7376_ _7376_/A _7376_/B _7376_/C vssd1 vssd1 vccd1 vccd1 _7378_/C sky130_fd_sc_hd__and3_1
XFILLER_103_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6327_ _6332_/B _6332_/C vssd1 vssd1 vccd1 vccd1 _6331_/A sky130_fd_sc_hd__nor2_1
X_4588_ _4588_/A vssd1 vssd1 vccd1 vccd1 _8582_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6258_ _6258_/A _6258_/B vssd1 vssd1 vccd1 vccd1 _6259_/B sky130_fd_sc_hd__xor2_1
X_5209_ _5233_/B _5209_/B _5209_/C _5223_/D vssd1 vssd1 vccd1 vccd1 _5210_/C sky130_fd_sc_hd__or4_1
X_6189_ _6187_/Y _6009_/B _6188_/Y vssd1 vssd1 vccd1 vccd1 _6230_/A sky130_fd_sc_hd__a21bo_2
XFILLER_84_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5560_ _5560_/A _5884_/B vssd1 vssd1 vccd1 vccd1 _5709_/A sky130_fd_sc_hd__or2_1
X_4511_ _4511_/A _4541_/B vssd1 vssd1 vccd1 vccd1 _4512_/A sky130_fd_sc_hd__or2_1
X_5491_ _5489_/X _5491_/B vssd1 vssd1 vccd1 vccd1 _5493_/B sky130_fd_sc_hd__and2b_1
X_4442_ _4443_/A vssd1 vssd1 vccd1 vccd1 _4442_/Y sky130_fd_sc_hd__inv_2
X_7230_ _7230_/A _7230_/B _7230_/C vssd1 vssd1 vccd1 vccd1 _7231_/A sky130_fd_sc_hd__nor3_1
XFILLER_104_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4373_ _4375_/A vssd1 vssd1 vccd1 vccd1 _4373_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7161_ _7159_/A _7159_/B _7160_/X vssd1 vssd1 vccd1 vccd1 _7291_/A sky130_fd_sc_hd__o21ba_1
X_7092_ _7101_/A _7101_/B _7093_/C vssd1 vssd1 vccd1 vccd1 _7105_/C sky130_fd_sc_hd__a21o_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6112_ _6111_/A _6111_/C _6117_/A vssd1 vssd1 vccd1 vccd1 _6113_/C sky130_fd_sc_hd__o21ai_1
X_6043_ _6043_/A _6043_/B vssd1 vssd1 vccd1 vccd1 _6044_/B sky130_fd_sc_hd__nand2_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7994_ _8076_/A _7994_/B vssd1 vssd1 vccd1 vccd1 _8078_/B sky130_fd_sc_hd__and2b_1
XFILLER_26_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6945_ _7096_/A _6945_/B vssd1 vssd1 vccd1 vccd1 _6945_/X sky130_fd_sc_hd__or2_1
XFILLER_26_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_2_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
X_6876_ _6876_/A _6876_/B vssd1 vssd1 vccd1 vccd1 _7349_/A sky130_fd_sc_hd__nor2_1
XFILLER_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8615_ _8733_/CLK _8615_/D vssd1 vssd1 vccd1 vccd1 _8615_/Q sky130_fd_sc_hd__dfxtp_2
X_5827_ _5827_/A _5827_/B vssd1 vssd1 vccd1 vccd1 _5828_/B sky130_fd_sc_hd__and2_1
X_8546_ _8547_/A _8560_/B vssd1 vssd1 vccd1 vccd1 _8548_/A sky130_fd_sc_hd__nor2_1
X_5758_ _6049_/A _6049_/B vssd1 vssd1 vccd1 vccd1 _5767_/A sky130_fd_sc_hd__and2_1
X_4709_ _5029_/A _5029_/B vssd1 vssd1 vccd1 vccd1 _4710_/A sky130_fd_sc_hd__nor2_1
X_8477_ _8477_/A _8477_/B vssd1 vssd1 vccd1 vccd1 _8478_/B sky130_fd_sc_hd__xnor2_1
X_7428_ _7428_/A _7428_/B vssd1 vssd1 vccd1 vccd1 _7462_/A sky130_fd_sc_hd__xnor2_1
X_5689_ _5692_/B _5692_/C vssd1 vssd1 vccd1 vccd1 _5690_/C sky130_fd_sc_hd__nand2_1
XFILLER_78_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7359_ _7455_/B _7447_/B _7359_/C vssd1 vssd1 vccd1 vccd1 _7362_/A sky130_fd_sc_hd__nand3_1
XFILLER_89_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6730_ _6730_/A _6730_/B vssd1 vssd1 vccd1 vccd1 _6829_/A sky130_fd_sc_hd__xnor2_1
X_4991_ _5196_/B _4991_/B _5169_/A vssd1 vssd1 vccd1 vccd1 _5164_/D sky130_fd_sc_hd__or3_1
XFILLER_51_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6661_ _6678_/A _6678_/B vssd1 vssd1 vccd1 vccd1 _6670_/B sky130_fd_sc_hd__xnor2_2
XFILLER_31_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6592_ _6592_/A _6592_/B vssd1 vssd1 vccd1 vccd1 _7501_/A sky130_fd_sc_hd__xnor2_1
XFILLER_31_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8400_ _8450_/A _8400_/B vssd1 vssd1 vccd1 vccd1 _8401_/B sky130_fd_sc_hd__nor2_1
X_5612_ _8662_/Q _7737_/B vssd1 vssd1 vccd1 vccd1 _5621_/B sky130_fd_sc_hd__and2b_1
X_5543_ _5560_/A _5992_/B vssd1 vssd1 vccd1 vccd1 _5574_/A sky130_fd_sc_hd__nor2_2
X_8331_ _8331_/A _8338_/A vssd1 vssd1 vccd1 vccd1 _8332_/B sky130_fd_sc_hd__xor2_1
X_8262_ _8262_/A _8262_/B vssd1 vssd1 vccd1 vccd1 _8430_/B sky130_fd_sc_hd__xnor2_2
X_5474_ _5474_/A _5503_/A vssd1 vssd1 vccd1 vccd1 _5499_/A sky130_fd_sc_hd__nand2_1
X_7213_ _6711_/A _7213_/B _7254_/C _7213_/D vssd1 vssd1 vccd1 vccd1 _7220_/B sky130_fd_sc_hd__and4b_1
X_4425_ _4425_/A vssd1 vssd1 vccd1 vccd1 _4425_/Y sky130_fd_sc_hd__inv_2
X_8193_ _8163_/A _8163_/B _8192_/Y vssd1 vssd1 vccd1 vccd1 _8274_/A sky130_fd_sc_hd__a21oi_2
XFILLER_98_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4356_ _4357_/A vssd1 vssd1 vccd1 vccd1 _4356_/Y sky130_fd_sc_hd__inv_2
X_7144_ _7154_/C _7154_/B _7185_/A vssd1 vssd1 vccd1 vccd1 _7190_/B sky130_fd_sc_hd__a21boi_1
XFILLER_58_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7075_ _7075_/A _7128_/B _7130_/B vssd1 vssd1 vccd1 vccd1 _7078_/A sky130_fd_sc_hd__or3_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6026_ _6026_/A _6026_/B vssd1 vssd1 vccd1 vccd1 _6043_/A sky130_fd_sc_hd__xnor2_1
XFILLER_104_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7977_ _8024_/A _7976_/B _7976_/C vssd1 vssd1 vccd1 vccd1 _7978_/C sky130_fd_sc_hd__a21o_1
X_6928_ _7054_/B _7430_/B _7007_/B vssd1 vssd1 vccd1 vccd1 _6934_/A sky130_fd_sc_hd__or3_1
XFILLER_42_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6859_ _6859_/A _6859_/B vssd1 vssd1 vccd1 vccd1 _6861_/B sky130_fd_sc_hd__xnor2_1
XFILLER_80_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8529_ _8529_/A _8529_/B vssd1 vssd1 vccd1 vccd1 _8529_/Y sky130_fd_sc_hd__nand2_1
XFILLER_89_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5190_ _5190_/A _5190_/B _5190_/C vssd1 vssd1 vccd1 vccd1 _5190_/X sky130_fd_sc_hd__or3_1
XFILLER_68_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7900_ _7945_/B _7945_/C _7945_/A vssd1 vssd1 vccd1 vccd1 _7928_/B sky130_fd_sc_hd__a21o_1
X_8880_ _8880_/A _4392_/Y vssd1 vssd1 vccd1 vccd1 io_out[17] sky130_fd_sc_hd__ebufn_8
XFILLER_48_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7831_ _7831_/A _7831_/B _7831_/C vssd1 vssd1 vccd1 vccd1 _7832_/B sky130_fd_sc_hd__or3_1
X_4974_ _5222_/A vssd1 vssd1 vccd1 vccd1 _5194_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_63_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7762_ _8399_/A _8122_/C _8122_/B _7761_/Y vssd1 vssd1 vccd1 vccd1 _7763_/B sky130_fd_sc_hd__o211a_1
X_6713_ _7409_/A _6713_/B vssd1 vssd1 vccd1 vccd1 _6768_/B sky130_fd_sc_hd__xnor2_1
X_7693_ _7759_/A _7759_/B vssd1 vssd1 vccd1 vccd1 _8118_/A sky130_fd_sc_hd__xor2_2
XFILLER_32_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6644_ _6759_/A vssd1 vssd1 vccd1 vccd1 _6797_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6575_ _6699_/A _7254_/B vssd1 vssd1 vccd1 vccd1 _6893_/C sky130_fd_sc_hd__nand2_1
X_8314_ _8314_/A _8314_/B vssd1 vssd1 vccd1 vccd1 _8386_/B sky130_fd_sc_hd__xnor2_2
X_5526_ _5873_/A _5992_/A vssd1 vssd1 vccd1 vccd1 _5532_/A sky130_fd_sc_hd__nor2_1
X_5457_ _6353_/A _4720_/A _6557_/B _6346_/A vssd1 vssd1 vccd1 vccd1 _5457_/X sky130_fd_sc_hd__o211a_1
X_8245_ _8489_/A _8279_/B vssd1 vssd1 vccd1 vccd1 _8246_/B sky130_fd_sc_hd__xor2_1
XFILLER_59_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4408_ _4432_/A vssd1 vssd1 vccd1 vccd1 _4413_/A sky130_fd_sc_hd__buf_6
XFILLER_99_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5388_ _5426_/A _5432_/A _5387_/X _8663_/Q vssd1 vssd1 vccd1 vccd1 _5389_/B sky130_fd_sc_hd__a31o_1
X_8176_ _8258_/B _8176_/B vssd1 vssd1 vccd1 vccd1 _8178_/B sky130_fd_sc_hd__xnor2_1
XFILLER_86_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7127_ _7127_/A _7127_/B vssd1 vssd1 vccd1 vccd1 _7143_/A sky130_fd_sc_hd__xnor2_1
X_4339_ _4464_/A vssd1 vssd1 vccd1 vccd1 _4344_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_101_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7058_ _7063_/B _7165_/B vssd1 vssd1 vccd1 vccd1 _7068_/A sky130_fd_sc_hd__xor2_1
XFILLER_59_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6009_ _6187_/A _6009_/B vssd1 vssd1 vccd1 vccd1 _6165_/B sky130_fd_sc_hd__xnor2_1
XFILLER_46_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4690_ _4690_/A vssd1 vssd1 vccd1 vccd1 _8603_/D sky130_fd_sc_hd__clkbuf_1
X_6360_ _6360_/A _6368_/B vssd1 vssd1 vccd1 vccd1 _6361_/B sky130_fd_sc_hd__or2b_1
X_5311_ _5323_/A vssd1 vssd1 vccd1 vccd1 _5311_/X sky130_fd_sc_hd__clkbuf_2
X_6291_ _6291_/A _6291_/B vssd1 vssd1 vccd1 vccd1 _6291_/Y sky130_fd_sc_hd__nor2_1
X_8030_ _8123_/S _8030_/B vssd1 vssd1 vccd1 vccd1 _8116_/A sky130_fd_sc_hd__xnor2_2
XFILLER_102_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5242_ _5236_/X _5237_/Y _5239_/X _5241_/X vssd1 vssd1 vccd1 vccd1 _5242_/X sky130_fd_sc_hd__o31a_1
X_5173_ _5173_/A _5173_/B vssd1 vssd1 vccd1 vccd1 _5173_/Y sky130_fd_sc_hd__nand2_1
Xinput1 active vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_6
XFILLER_96_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8932_ _8932_/A _4453_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[31] sky130_fd_sc_hd__ebufn_8
X_8863_ _8863_/A _4462_/Y vssd1 vssd1 vccd1 vccd1 io_out[0] sky130_fd_sc_hd__ebufn_8
XFILLER_83_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7814_ _7903_/C _7814_/B vssd1 vssd1 vccd1 vccd1 _7815_/B sky130_fd_sc_hd__xor2_1
XFILLER_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4957_ _4957_/A _5175_/B vssd1 vssd1 vccd1 vccd1 _4958_/B sky130_fd_sc_hd__and2_1
XFILLER_51_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7745_ _7835_/A _8145_/A vssd1 vssd1 vccd1 vccd1 _7813_/B sky130_fd_sc_hd__nor2_2
X_4888_ _4996_/A _5099_/A vssd1 vssd1 vccd1 vccd1 _5038_/A sky130_fd_sc_hd__or2_2
X_7676_ _8733_/Q _7677_/B vssd1 vssd1 vccd1 vccd1 _7769_/A sky130_fd_sc_hd__nor2_2
X_6627_ _6663_/A vssd1 vssd1 vccd1 vccd1 _6688_/A sky130_fd_sc_hd__clkbuf_2
X_6558_ _6558_/A _6558_/B vssd1 vssd1 vccd1 vccd1 _6559_/B sky130_fd_sc_hd__nor2_2
XFILLER_20_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6489_ _8699_/Q vssd1 vssd1 vccd1 vccd1 _6509_/A sky130_fd_sc_hd__clkbuf_2
X_5509_ _5567_/B _5896_/A _5509_/C vssd1 vssd1 vccd1 vccd1 _6019_/B sky130_fd_sc_hd__and3_1
X_8228_ _8228_/A _8338_/B vssd1 vssd1 vccd1 vccd1 _8231_/A sky130_fd_sc_hd__xnor2_1
X_8159_ _8256_/A _8159_/B vssd1 vssd1 vccd1 vccd1 _8161_/B sky130_fd_sc_hd__nor2_1
XFILLER_87_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5860_ _6119_/A _5941_/C _5953_/A vssd1 vssd1 vccd1 vccd1 _6196_/A sky130_fd_sc_hd__o21a_2
XFILLER_46_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4811_ _4828_/A _4847_/A _4818_/B vssd1 vssd1 vccd1 vccd1 _4830_/A sky130_fd_sc_hd__or3_2
XFILLER_61_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5791_ _5881_/B _5882_/B vssd1 vssd1 vccd1 vccd1 _5800_/A sky130_fd_sc_hd__xnor2_1
X_7530_ _7526_/A _5308_/X _6508_/A _7529_/Y vssd1 vssd1 vccd1 vccd1 _8712_/D sky130_fd_sc_hd__a22o_1
X_4742_ _8613_/Q vssd1 vssd1 vccd1 vccd1 _4848_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_14_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7461_ _7461_/A _7461_/B vssd1 vssd1 vccd1 vccd1 _7462_/B sky130_fd_sc_hd__xnor2_2
X_4673_ _4661_/A _4763_/A _4702_/B _4672_/X vssd1 vssd1 vccd1 vccd1 _8602_/D sky130_fd_sc_hd__o211a_1
X_6412_ _8678_/Q _6413_/B vssd1 vssd1 vccd1 vccd1 _6418_/C sky130_fd_sc_hd__and2_1
X_7392_ _7392_/A _7399_/A vssd1 vssd1 vccd1 vccd1 _7397_/A sky130_fd_sc_hd__xnor2_1
X_6343_ _8668_/Q _6343_/B vssd1 vssd1 vccd1 vccd1 _6343_/Y sky130_fd_sc_hd__xnor2_1
X_6274_ _6274_/A _6274_/B vssd1 vssd1 vccd1 vccd1 _6275_/B sky130_fd_sc_hd__xor2_1
X_5225_ _5120_/A _5199_/C _5222_/X _5224_/X vssd1 vssd1 vccd1 vccd1 _5226_/D sky130_fd_sc_hd__o31a_1
X_8013_ _7936_/A _7938_/A _8021_/B _8012_/X vssd1 vssd1 vccd1 vccd1 _8019_/A sky130_fd_sc_hd__o211a_1
XFILLER_69_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5156_ _5154_/X _5155_/X _4916_/A vssd1 vssd1 vccd1 vccd1 _5156_/X sky130_fd_sc_hd__a21o_1
XFILLER_56_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5087_ _5087_/A _5087_/B vssd1 vssd1 vccd1 vccd1 _5119_/A sky130_fd_sc_hd__and2_1
XFILLER_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8915_ _8915_/A _4433_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[14] sky130_fd_sc_hd__ebufn_8
XFILLER_44_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8846_ _8846_/A _4351_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[15] sky130_fd_sc_hd__ebufn_8
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5989_ _5989_/A _5989_/B vssd1 vssd1 vccd1 vccd1 _6200_/A sky130_fd_sc_hd__xnor2_1
XFILLER_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7728_ _7728_/A vssd1 vssd1 vccd1 vccd1 _8206_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_20_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7659_ _7835_/B vssd1 vssd1 vccd1 vccd1 _8281_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_21_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_3_4_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_9_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5010_ _5028_/B _4992_/X _5005_/X _5009_/X vssd1 vssd1 vccd1 vccd1 _5010_/X sky130_fd_sc_hd__o211a_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6961_ _6960_/B _6960_/C _7348_/C vssd1 vssd1 vccd1 vccd1 _6962_/C sky130_fd_sc_hd__a21oi_1
XFILLER_66_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8700_ _8733_/CLK _8700_/D vssd1 vssd1 vccd1 vccd1 _8700_/Q sky130_fd_sc_hd__dfxtp_1
X_6892_ _6892_/A _6892_/B vssd1 vssd1 vccd1 vccd1 _6954_/A sky130_fd_sc_hd__xor2_1
X_5912_ _6238_/A _5938_/B vssd1 vssd1 vccd1 vccd1 _5913_/B sky130_fd_sc_hd__xnor2_1
XFILLER_46_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8631_ _8734_/CLK _8631_/D vssd1 vssd1 vccd1 vccd1 _8631_/Q sky130_fd_sc_hd__dfxtp_1
X_5843_ _5924_/B _5843_/B vssd1 vssd1 vccd1 vccd1 _5845_/B sky130_fd_sc_hd__xnor2_1
XFILLER_34_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8780__47 vssd1 vssd1 vccd1 vccd1 _8780__47/HI _8889_/A sky130_fd_sc_hd__conb_1
X_8562_ _8554_/B _8562_/B vssd1 vssd1 vccd1 vccd1 _8563_/C sky130_fd_sc_hd__and2b_1
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7513_ _7513_/A vssd1 vssd1 vccd1 vccd1 _8709_/D sky130_fd_sc_hd__clkbuf_1
X_5774_ _5726_/A _5726_/B _5721_/A _5721_/B vssd1 vssd1 vccd1 vccd1 _5856_/A sky130_fd_sc_hd__o2bb2a_1
X_4725_ _4801_/B _4726_/B vssd1 vssd1 vccd1 vccd1 _4727_/B sky130_fd_sc_hd__or2_1
X_8493_ _8493_/A _8493_/B _8493_/C vssd1 vssd1 vccd1 vccd1 _8512_/A sky130_fd_sc_hd__and3_1
X_7444_ _7444_/A _7444_/B vssd1 vssd1 vccd1 vccd1 _7445_/B sky130_fd_sc_hd__xnor2_1
X_4656_ _5154_/A vssd1 vssd1 vccd1 vccd1 _5153_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7375_ _6985_/A _6985_/B _6985_/C _6984_/B _6984_/A vssd1 vssd1 vccd1 vccd1 _7376_/C
+ sky130_fd_sc_hd__a32o_1
X_4587_ _4587_/A _4612_/B _4587_/C vssd1 vssd1 vccd1 vccd1 _4588_/A sky130_fd_sc_hd__and3_1
X_6326_ _6319_/X _6324_/X _6325_/X _8664_/Q vssd1 vssd1 vccd1 vccd1 _8664_/D sky130_fd_sc_hd__o2bb2a_1
XFILLER_88_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6257_ _6219_/S _6220_/A _6256_/X vssd1 vssd1 vccd1 vccd1 _6258_/B sky130_fd_sc_hd__a21bo_1
XFILLER_88_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5208_ _5208_/A _5224_/B _5208_/C _5208_/D vssd1 vssd1 vccd1 vccd1 _5208_/X sky130_fd_sc_hd__or4_1
X_6188_ _6188_/A _6188_/B vssd1 vssd1 vccd1 vccd1 _6188_/Y sky130_fd_sc_hd__nand2_1
X_5139_ _5223_/A _5202_/C _5139_/C _5139_/D vssd1 vssd1 vccd1 vccd1 _5139_/X sky130_fd_sc_hd__or4_1
XFILLER_57_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4510_ _4660_/A _4790_/A _4820_/B _4787_/A vssd1 vssd1 vccd1 vccd1 _4541_/B sky130_fd_sc_hd__a31oi_2
X_5490_ _8611_/Q _8674_/Q vssd1 vssd1 vccd1 vccd1 _5491_/B sky130_fd_sc_hd__or2b_1
X_4441_ _4443_/A vssd1 vssd1 vccd1 vccd1 _4441_/Y sky130_fd_sc_hd__inv_2
X_7160_ _7195_/A _7195_/B vssd1 vssd1 vccd1 vccd1 _7160_/X sky130_fd_sc_hd__and2b_1
X_4372_ _4375_/A vssd1 vssd1 vccd1 vccd1 _4372_/Y sky130_fd_sc_hd__inv_2
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6111_ _6111_/A _6117_/A _6111_/C vssd1 vssd1 vccd1 vccd1 _6143_/A sky130_fd_sc_hd__or3_2
X_7091_ _7091_/A _7091_/B vssd1 vssd1 vccd1 vccd1 _7093_/C sky130_fd_sc_hd__xor2_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6042_ _6043_/A _6043_/B vssd1 vssd1 vccd1 vccd1 _6051_/A sky130_fd_sc_hd__or2_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8825__92 vssd1 vssd1 vccd1 vccd1 _8825__92/HI _8934_/A sky130_fd_sc_hd__conb_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7993_ _8008_/A _7993_/B _7998_/A vssd1 vssd1 vccd1 vccd1 _7994_/B sky130_fd_sc_hd__or3b_1
XFILLER_26_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6944_ _6944_/A _6944_/B vssd1 vssd1 vccd1 vccd1 _7119_/B sky130_fd_sc_hd__xnor2_1
XFILLER_81_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6875_ _7364_/B _7355_/A vssd1 vssd1 vccd1 vccd1 _6882_/A sky130_fd_sc_hd__nor2_1
X_8614_ _8671_/CLK _8614_/D vssd1 vssd1 vccd1 vccd1 _8614_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5826_ _5827_/A _5827_/B vssd1 vssd1 vccd1 vccd1 _5922_/B sky130_fd_sc_hd__nor2_1
X_5757_ _5757_/A _5770_/B vssd1 vssd1 vccd1 vccd1 _6018_/A sky130_fd_sc_hd__xnor2_1
XFILLER_22_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8545_ _8545_/A vssd1 vssd1 vccd1 vccd1 _8730_/D sky130_fd_sc_hd__clkbuf_1
X_4708_ _6553_/B _5080_/B vssd1 vssd1 vccd1 vccd1 _5029_/B sky130_fd_sc_hd__nor2_1
X_8476_ _8476_/A _8476_/B vssd1 vssd1 vccd1 vccd1 _8477_/B sky130_fd_sc_hd__xnor2_1
X_7427_ _7427_/A _7427_/B vssd1 vssd1 vccd1 vccd1 _7428_/B sky130_fd_sc_hd__xnor2_1
X_5688_ _6026_/A _6026_/B vssd1 vssd1 vccd1 vccd1 _5692_/C sky130_fd_sc_hd__or2_1
X_4639_ _4643_/C _4645_/B _4639_/C vssd1 vssd1 vccd1 vccd1 _4640_/A sky130_fd_sc_hd__and3b_1
X_7358_ _6978_/B _6978_/C _6978_/A vssd1 vssd1 vccd1 vccd1 _7359_/C sky130_fd_sc_hd__a21bo_1
XFILLER_89_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7289_ _7289_/A _7250_/A vssd1 vssd1 vccd1 vccd1 _7478_/A sky130_fd_sc_hd__or2b_1
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6309_ _6309_/A _6309_/B vssd1 vssd1 vccd1 vccd1 _6309_/Y sky130_fd_sc_hd__nor2_1
XFILLER_103_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4990_ _4990_/A _4990_/B vssd1 vssd1 vccd1 vccd1 _5245_/D sky130_fd_sc_hd__nor2_2
XFILLER_16_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6660_ _6579_/A _6579_/B _6631_/A vssd1 vssd1 vccd1 vccd1 _6678_/B sky130_fd_sc_hd__a21boi_2
X_8750__17 vssd1 vssd1 vccd1 vccd1 _8750__17/HI _8845_/A sky130_fd_sc_hd__conb_1
X_6591_ _7454_/A _6578_/B _6807_/A vssd1 vssd1 vccd1 vccd1 _6592_/B sky130_fd_sc_hd__o21a_1
X_5611_ _5660_/A _5661_/A _5661_/B _5599_/X _5603_/A vssd1 vssd1 vccd1 vccd1 _5619_/B
+ sky130_fd_sc_hd__a311o_1
X_5542_ _5884_/B vssd1 vssd1 vccd1 vccd1 _5992_/B sky130_fd_sc_hd__clkbuf_2
X_8330_ _8330_/A _8450_/A vssd1 vssd1 vccd1 vccd1 _8338_/A sky130_fd_sc_hd__nor2_1
X_8261_ _8271_/A _8271_/B vssd1 vssd1 vccd1 vccd1 _8262_/B sky130_fd_sc_hd__xor2_2
X_5473_ _5519_/A _5519_/B vssd1 vssd1 vccd1 vccd1 _5503_/A sky130_fd_sc_hd__xor2_2
X_7212_ _7212_/A _7212_/B vssd1 vssd1 vccd1 vccd1 _7220_/A sky130_fd_sc_hd__xor2_1
X_8192_ _8192_/A _8192_/B vssd1 vssd1 vccd1 vccd1 _8192_/Y sky130_fd_sc_hd__nor2_1
X_4424_ _4425_/A vssd1 vssd1 vccd1 vccd1 _4424_/Y sky130_fd_sc_hd__inv_2
X_4355_ _4357_/A vssd1 vssd1 vccd1 vccd1 _4355_/Y sky130_fd_sc_hd__inv_2
X_7143_ _7143_/A _7143_/B _7143_/C vssd1 vssd1 vccd1 vccd1 _7185_/A sky130_fd_sc_hd__nand3_1
XFILLER_98_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7074_ _7082_/A _7074_/B _7074_/C vssd1 vssd1 vccd1 vccd1 _7130_/B sky130_fd_sc_hd__or3_2
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6025_ _6024_/A _6024_/C _6024_/B vssd1 vssd1 vccd1 vccd1 _6045_/B sky130_fd_sc_hd__a21oi_1
XFILLER_39_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7976_ _8024_/A _7976_/B _7976_/C vssd1 vssd1 vccd1 vccd1 _8024_/B sky130_fd_sc_hd__nand3_1
XFILLER_14_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6927_ _6927_/A vssd1 vssd1 vccd1 vccd1 _7430_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6858_ _6914_/B _6857_/Y _7409_/B vssd1 vssd1 vccd1 vccd1 _6859_/B sky130_fd_sc_hd__a21oi_1
XFILLER_50_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5809_ _5856_/A _5856_/B vssd1 vssd1 vccd1 vccd1 _5829_/A sky130_fd_sc_hd__xor2_2
XFILLER_22_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6789_ _6789_/A _6789_/B _6789_/C vssd1 vssd1 vccd1 vccd1 _6790_/B sky130_fd_sc_hd__and3_1
XFILLER_13_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8528_ _8529_/A _8529_/B vssd1 vssd1 vccd1 vccd1 _8533_/B sky130_fd_sc_hd__or2_1
X_8459_ _8459_/A _8459_/B vssd1 vssd1 vccd1 vccd1 _8463_/A sky130_fd_sc_hd__xnor2_1
XFILLER_2_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7830_ _7831_/B _7831_/C _7831_/A vssd1 vssd1 vccd1 vccd1 _8101_/A sky130_fd_sc_hd__o21ai_2
XFILLER_91_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4973_ _5056_/A _4973_/B vssd1 vssd1 vccd1 vccd1 _4973_/X sky130_fd_sc_hd__or2_1
XFILLER_51_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7761_ _7862_/A _8130_/A vssd1 vssd1 vccd1 vccd1 _7761_/Y sky130_fd_sc_hd__nand2_1
X_6712_ _6708_/X _7369_/A _6785_/A vssd1 vssd1 vccd1 vccd1 _6713_/B sky130_fd_sc_hd__a21oi_2
X_7692_ _7712_/A _7712_/B _7713_/B _7691_/X _7689_/A vssd1 vssd1 vccd1 vccd1 _7759_/B
+ sky130_fd_sc_hd__a311o_4
X_6643_ _7102_/A _7370_/A vssd1 vssd1 vccd1 vccd1 _7103_/A sky130_fd_sc_hd__nor2_2
XFILLER_32_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6574_ _6735_/A vssd1 vssd1 vccd1 vccd1 _7254_/B sky130_fd_sc_hd__clkbuf_2
X_8313_ _8289_/A _8489_/B _8312_/Y vssd1 vssd1 vccd1 vccd1 _8314_/B sky130_fd_sc_hd__o21ba_1
X_5525_ _5525_/A vssd1 vssd1 vccd1 vccd1 _5992_/A sky130_fd_sc_hd__clkbuf_2
X_8244_ _8370_/A _8147_/X _8196_/X vssd1 vssd1 vccd1 vccd1 _8279_/B sky130_fd_sc_hd__o21a_1
X_5456_ _5456_/A vssd1 vssd1 vccd1 vccd1 _6346_/A sky130_fd_sc_hd__inv_2
X_4407_ input1/X vssd1 vssd1 vccd1 vccd1 _4432_/A sky130_fd_sc_hd__clkbuf_2
X_8175_ _8087_/A _8087_/C _8087_/B vssd1 vssd1 vccd1 vccd1 _8176_/B sky130_fd_sc_hd__a21boi_1
X_5387_ _5400_/A _8657_/Q _5411_/B _5404_/B vssd1 vssd1 vccd1 vccd1 _5387_/X sky130_fd_sc_hd__a211o_1
XFILLER_101_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7126_ _7125_/A _7125_/B _7125_/C _7125_/D vssd1 vssd1 vccd1 vccd1 _7154_/B sky130_fd_sc_hd__o22ai_1
X_4338_ _4338_/A vssd1 vssd1 vccd1 vccd1 _4338_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7057_ _7146_/A _7057_/B vssd1 vssd1 vccd1 vccd1 _7151_/A sky130_fd_sc_hd__xnor2_2
XFILLER_74_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6008_ _6188_/A _6188_/B vssd1 vssd1 vccd1 vccd1 _6009_/B sky130_fd_sc_hd__xor2_1
XFILLER_27_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7959_ _8026_/B _7958_/C _7958_/A vssd1 vssd1 vccd1 vccd1 _7966_/B sky130_fd_sc_hd__a21o_1
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5310_ _5314_/C _5310_/B vssd1 vssd1 vccd1 vccd1 _8637_/D sky130_fd_sc_hd__nor2_1
X_6290_ _6290_/A _6290_/B vssd1 vssd1 vccd1 vccd1 _6293_/A sky130_fd_sc_hd__xnor2_4
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5241_ _4923_/A _5132_/C _5127_/D _5240_/X _5067_/C vssd1 vssd1 vccd1 vccd1 _5241_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_96_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5172_ _5172_/A _5172_/B _5240_/D _5175_/D vssd1 vssd1 vccd1 vccd1 _5172_/X sky130_fd_sc_hd__or4_1
XFILLER_96_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput2 io_in[10] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__buf_4
X_8931_ _8931_/A _4452_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[30] sky130_fd_sc_hd__ebufn_8
XFILLER_68_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8862_ _8862_/A _4371_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[31] sky130_fd_sc_hd__ebufn_8
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7813_ _7813_/A _7813_/B vssd1 vssd1 vccd1 vccd1 _7814_/B sky130_fd_sc_hd__xnor2_1
XFILLER_51_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7744_ _8515_/A _8304_/A vssd1 vssd1 vccd1 vccd1 _7748_/A sky130_fd_sc_hd__nor2_1
X_4956_ _4956_/A vssd1 vssd1 vccd1 vccd1 _5175_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_51_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4887_ _5107_/A _4964_/B _5111_/B vssd1 vssd1 vccd1 vccd1 _5099_/A sky130_fd_sc_hd__or3_1
X_7675_ _7675_/A _7675_/B vssd1 vssd1 vccd1 vccd1 _7750_/A sky130_fd_sc_hd__xnor2_1
X_6626_ _8620_/Q _6536_/A vssd1 vssd1 vccd1 vccd1 _6663_/A sky130_fd_sc_hd__or2b_1
X_6557_ _8711_/Q _6557_/B vssd1 vssd1 vccd1 vccd1 _6558_/B sky130_fd_sc_hd__and2b_1
X_5508_ _5872_/B _5993_/A vssd1 vssd1 vccd1 vccd1 _5509_/C sky130_fd_sc_hd__or2_1
X_6488_ _8700_/Q vssd1 vssd1 vccd1 vccd1 _6515_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5439_ _5439_/A vssd1 vssd1 vccd1 vccd1 _5540_/A sky130_fd_sc_hd__clkbuf_2
X_8227_ _7885_/A _8204_/A _8410_/A _8220_/B vssd1 vssd1 vccd1 vccd1 _8338_/B sky130_fd_sc_hd__o22a_1
X_8158_ _8158_/A _8158_/B vssd1 vssd1 vccd1 vccd1 _8159_/B sky130_fd_sc_hd__nor2_1
XFILLER_87_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7109_ _7109_/A _7109_/B vssd1 vssd1 vccd1 vccd1 _7113_/B sky130_fd_sc_hd__xnor2_1
XFILLER_59_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8089_ _8258_/A _8089_/B vssd1 vssd1 vccd1 vccd1 _8091_/B sky130_fd_sc_hd__nor2_1
XFILLER_74_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8786__53 vssd1 vssd1 vccd1 vccd1 _8786__53/HI _8895_/A sky130_fd_sc_hd__conb_1
XFILLER_27_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_6_0_wb_clk_i clkbuf_4_7_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _8733_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_27_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4810_ _4848_/B _4848_/C vssd1 vssd1 vccd1 vccd1 _4818_/B sky130_fd_sc_hd__nand2_1
XFILLER_21_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5790_ _5790_/A _5790_/B vssd1 vssd1 vccd1 vccd1 _5882_/B sky130_fd_sc_hd__xnor2_1
X_4741_ _4891_/A _4752_/A _4740_/X vssd1 vssd1 vccd1 vccd1 _8612_/D sky130_fd_sc_hd__a21oi_1
X_7460_ _7460_/A _7460_/B vssd1 vssd1 vccd1 vccd1 _7461_/B sky130_fd_sc_hd__xnor2_1
X_4672_ _4727_/A vssd1 vssd1 vccd1 vccd1 _4672_/X sky130_fd_sc_hd__clkbuf_2
X_6411_ _6411_/A vssd1 vssd1 vccd1 vccd1 _8677_/D sky130_fd_sc_hd__clkbuf_1
X_7391_ _7391_/A _7391_/B vssd1 vssd1 vccd1 vccd1 _7399_/A sky130_fd_sc_hd__xnor2_1
X_6342_ _6342_/A _6342_/B vssd1 vssd1 vccd1 vccd1 _6343_/B sky130_fd_sc_hd__nand2_1
X_6273_ _6194_/A _5973_/A _6273_/S vssd1 vssd1 vccd1 vccd1 _6274_/B sky130_fd_sc_hd__mux2_1
XFILLER_88_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5224_ _5231_/B _5224_/B _5224_/C vssd1 vssd1 vccd1 vccd1 _5224_/X sky130_fd_sc_hd__or3_1
X_8012_ _8021_/A _8011_/B _8011_/C vssd1 vssd1 vccd1 vccd1 _8012_/X sky130_fd_sc_hd__a21o_1
XFILLER_84_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5155_ _5155_/A _5155_/B _5155_/C vssd1 vssd1 vccd1 vccd1 _5155_/X sky130_fd_sc_hd__or3_1
XFILLER_56_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5086_ _5227_/A _5086_/B vssd1 vssd1 vccd1 vccd1 _5109_/D sky130_fd_sc_hd__or2_1
XFILLER_84_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8914_ _8914_/A _4430_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[13] sky130_fd_sc_hd__ebufn_8
X_8845_ _8845_/A _4350_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[14] sky130_fd_sc_hd__ebufn_8
XFILLER_24_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5988_ _6191_/A _6191_/B vssd1 vssd1 vccd1 vccd1 _5989_/B sky130_fd_sc_hd__xor2_1
X_4939_ _4979_/A _5207_/B _5245_/B _5192_/D vssd1 vssd1 vccd1 vccd1 _4939_/X sky130_fd_sc_hd__or4_1
XFILLER_12_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7727_ _7833_/A _7727_/B vssd1 vssd1 vccd1 vccd1 _7841_/A sky130_fd_sc_hd__nand2_1
X_7658_ _7722_/A _7666_/B vssd1 vssd1 vccd1 vccd1 _7835_/B sky130_fd_sc_hd__xnor2_2
X_6609_ _7280_/A _6617_/A vssd1 vssd1 vccd1 vccd1 _6914_/A sky130_fd_sc_hd__nand2_4
XFILLER_20_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7589_ _8717_/Q _7590_/A vssd1 vssd1 vccd1 vccd1 _7591_/A sky130_fd_sc_hd__or2b_1
XFILLER_94_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6960_ _7348_/C _6960_/B _6960_/C vssd1 vssd1 vccd1 vccd1 _7361_/A sky130_fd_sc_hd__and3_1
XFILLER_81_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5911_ _6174_/A _5816_/B _5862_/Y vssd1 vssd1 vccd1 vccd1 _5938_/B sky130_fd_sc_hd__o21ai_1
X_6891_ _6958_/A vssd1 vssd1 vccd1 vccd1 _6892_/B sky130_fd_sc_hd__clkbuf_2
X_8630_ _8734_/CLK _8630_/D vssd1 vssd1 vccd1 vccd1 _8630_/Q sky130_fd_sc_hd__dfxtp_1
X_5842_ _5842_/A _5924_/A vssd1 vssd1 vccd1 vccd1 _5843_/B sky130_fd_sc_hd__nor2_1
X_8561_ _8569_/A _8561_/B vssd1 vssd1 vccd1 vccd1 _8563_/B sky130_fd_sc_hd__or2_1
X_5773_ _5756_/A _5756_/B _5772_/X vssd1 vssd1 vccd1 vccd1 _5830_/A sky130_fd_sc_hd__a21oi_1
XFILLER_21_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7512_ _5362_/A _6507_/A _7516_/A vssd1 vssd1 vccd1 vccd1 _7513_/A sky130_fd_sc_hd__mux2_1
X_4724_ _4724_/A vssd1 vssd1 vccd1 vccd1 _8608_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8492_ _8492_/A _8492_/B vssd1 vssd1 vccd1 vccd1 _8493_/C sky130_fd_sc_hd__xnor2_1
X_7443_ _7443_/A _7443_/B vssd1 vssd1 vccd1 vccd1 _7444_/B sky130_fd_sc_hd__xnor2_1
X_4655_ _4923_/A vssd1 vssd1 vccd1 vccd1 _5154_/A sky130_fd_sc_hd__clkbuf_2
X_7374_ _7447_/D _7373_/B _7373_/C vssd1 vssd1 vccd1 vccd1 _7376_/B sky130_fd_sc_hd__a21o_1
X_4586_ _8582_/Q _8581_/Q vssd1 vssd1 vccd1 vccd1 _4587_/C sky130_fd_sc_hd__nand2_1
X_6325_ _7537_/B vssd1 vssd1 vccd1 vccd1 _6325_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_103_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6256_ _6204_/A _5987_/A _6219_/S _6220_/A _6220_/B vssd1 vssd1 vccd1 vccd1 _6256_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_88_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5207_ _5207_/A _5207_/B _5231_/A _5207_/D vssd1 vssd1 vccd1 vccd1 _5208_/D sky130_fd_sc_hd__or4_1
XFILLER_69_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6187_ _6187_/A vssd1 vssd1 vccd1 vccd1 _6187_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5138_ _5138_/A vssd1 vssd1 vccd1 vccd1 _5223_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5069_ _5175_/A _5087_/A _5087_/B _5130_/A vssd1 vssd1 vccd1 vccd1 _5069_/X sky130_fd_sc_hd__a31o_1
X_8756__23 vssd1 vssd1 vccd1 vccd1 _8756__23/HI _8851_/A sky130_fd_sc_hd__conb_1
XFILLER_72_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4440_ _4443_/A vssd1 vssd1 vccd1 vccd1 _4440_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4371_ _4375_/A vssd1 vssd1 vccd1 vccd1 _4371_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6110_ _6110_/A _6110_/B vssd1 vssd1 vccd1 vccd1 _6111_/C sky130_fd_sc_hd__and2_1
X_7090_ _7087_/X _7136_/B _7089_/Y vssd1 vssd1 vccd1 vccd1 _7101_/B sky130_fd_sc_hd__a21bo_2
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6041_ _5680_/A _6027_/X _6036_/B _6040_/Y vssd1 vssd1 vccd1 vccd1 _6043_/B sky130_fd_sc_hd__o31a_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7992_ _8008_/A _7993_/B _7998_/A vssd1 vssd1 vccd1 vccd1 _8076_/A sky130_fd_sc_hd__o21ba_1
X_6943_ _6944_/A _6944_/B vssd1 vssd1 vccd1 vccd1 _6943_/Y sky130_fd_sc_hd__nand2_1
X_6874_ _7213_/B _7355_/A _7352_/B vssd1 vssd1 vccd1 vccd1 _6883_/A sky130_fd_sc_hd__a21oi_2
XFILLER_34_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8613_ _8671_/CLK _8613_/D vssd1 vssd1 vccd1 vccd1 _8613_/Q sky130_fd_sc_hd__dfxtp_1
X_5825_ _5922_/A _5825_/B vssd1 vssd1 vccd1 vccd1 _5827_/B sky130_fd_sc_hd__or2_1
XFILLER_34_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5756_ _5756_/A _5756_/B vssd1 vssd1 vccd1 vccd1 _5770_/B sky130_fd_sc_hd__xor2_1
X_8544_ _8544_/A _8544_/B vssd1 vssd1 vccd1 vccd1 _8545_/A sky130_fd_sc_hd__and2_1
X_4707_ _4707_/A _5053_/A vssd1 vssd1 vccd1 vccd1 _5080_/B sky130_fd_sc_hd__nor2_2
X_8475_ _8368_/B _8311_/A _8368_/Y vssd1 vssd1 vccd1 vccd1 _8476_/B sky130_fd_sc_hd__a21oi_1
X_5687_ _5687_/A _5687_/B vssd1 vssd1 vccd1 vccd1 _6026_/B sky130_fd_sc_hd__xnor2_1
X_7426_ _7388_/A _7387_/B _7387_/A vssd1 vssd1 vccd1 vccd1 _7427_/B sky130_fd_sc_hd__o21ba_1
X_4638_ _8596_/Q _8597_/Q _4632_/B _8598_/Q vssd1 vssd1 vccd1 vccd1 _4639_/C sky130_fd_sc_hd__a31o_1
X_7357_ _7355_/B _7355_/C _7355_/A vssd1 vssd1 vccd1 vccd1 _7447_/B sky130_fd_sc_hd__o21ai_2
X_4569_ input2/X vssd1 vssd1 vccd1 vccd1 _7499_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7288_ _7230_/B _7230_/C _7230_/A vssd1 vssd1 vccd1 vccd1 _7479_/A sky130_fd_sc_hd__o21ai_1
XFILLER_1_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6308_ _6311_/A _6311_/B _6154_/X vssd1 vssd1 vccd1 vccd1 _6309_/B sky130_fd_sc_hd__a21oi_1
X_6239_ _6239_/A _6239_/B vssd1 vssd1 vccd1 vccd1 _6239_/Y sky130_fd_sc_hd__nand2_1
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6590_ _6590_/A _7009_/B vssd1 vssd1 vccd1 vccd1 _6807_/A sky130_fd_sc_hd__nor2_1
X_5610_ _7737_/B _8662_/Q vssd1 vssd1 vccd1 vccd1 _5610_/X sky130_fd_sc_hd__or2b_1
X_5541_ _5541_/A vssd1 vssd1 vccd1 vccd1 _5884_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_8_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8260_ _8260_/A _8260_/B vssd1 vssd1 vccd1 vccd1 _8271_/B sky130_fd_sc_hd__xnor2_2
X_7211_ _7211_/A _7069_/A vssd1 vssd1 vccd1 vccd1 _7215_/A sky130_fd_sc_hd__or2b_1
X_5472_ _5475_/A _5475_/B _5447_/A vssd1 vssd1 vccd1 vccd1 _5519_/B sky130_fd_sc_hd__a21oi_2
X_4423_ _4425_/A vssd1 vssd1 vccd1 vccd1 _4423_/Y sky130_fd_sc_hd__inv_2
X_8191_ _8181_/A _8181_/B _8190_/X vssd1 vssd1 vccd1 vccd1 _8271_/A sky130_fd_sc_hd__a21boi_2
X_4354_ _4357_/A vssd1 vssd1 vccd1 vccd1 _4354_/Y sky130_fd_sc_hd__inv_2
X_7142_ _7141_/B _7141_/C _7141_/A vssd1 vssd1 vccd1 vccd1 _7143_/C sky130_fd_sc_hd__a21o_1
X_7073_ _7148_/A _7072_/X _6842_/Y vssd1 vssd1 vccd1 vccd1 _7151_/B sky130_fd_sc_hd__o21a_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6024_ _6024_/A _6024_/B _6024_/C vssd1 vssd1 vccd1 vccd1 _6046_/A sky130_fd_sc_hd__and3_1
XFILLER_100_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7975_ _8046_/A _7975_/B vssd1 vssd1 vccd1 vccd1 _7976_/C sky130_fd_sc_hd__xnor2_1
X_6926_ _6926_/A _6926_/B vssd1 vssd1 vccd1 vccd1 _6935_/A sky130_fd_sc_hd__nor2_1
XFILLER_81_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6857_ _6857_/A _6857_/B vssd1 vssd1 vccd1 vccd1 _6857_/Y sky130_fd_sc_hd__nand2_1
XFILLER_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6788_ _6789_/A _6789_/B _6789_/C vssd1 vssd1 vccd1 vccd1 _6790_/A sky130_fd_sc_hd__a21oi_1
XFILLER_50_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5808_ _5808_/A _5808_/B vssd1 vssd1 vccd1 vccd1 _5856_/B sky130_fd_sc_hd__xnor2_1
X_5739_ _5742_/A _5739_/B vssd1 vssd1 vccd1 vccd1 _5945_/A sky130_fd_sc_hd__nand2_2
X_8527_ _4771_/X _8520_/X _8525_/X _8526_/Y vssd1 vssd1 vccd1 vccd1 _8726_/D sky130_fd_sc_hd__a31oi_1
XFILLER_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8458_ _8401_/A _8401_/B _8402_/B _8195_/A vssd1 vssd1 vccd1 vccd1 _8459_/B sky130_fd_sc_hd__a22o_1
X_7409_ _7409_/A _7409_/B vssd1 vssd1 vccd1 vccd1 _7409_/Y sky130_fd_sc_hd__nor2_1
X_8389_ _8473_/S _8310_/B _8312_/B vssd1 vssd1 vccd1 vccd1 _8460_/B sky130_fd_sc_hd__a21bo_1
XFILLER_89_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8810__77 vssd1 vssd1 vccd1 vccd1 _8810__77/HI _8919_/A sky130_fd_sc_hd__conb_1
XFILLER_51_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4972_ _4692_/A _4960_/B _4954_/X _4971_/X _4697_/X vssd1 vssd1 vccd1 vccd1 _4973_/B
+ sky130_fd_sc_hd__o32a_1
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7760_ _7862_/A vssd1 vssd1 vccd1 vccd1 _8399_/A sky130_fd_sc_hd__buf_2
X_6711_ _6711_/A _7370_/A vssd1 vssd1 vccd1 vccd1 _6785_/A sky130_fd_sc_hd__nor2_1
X_7691_ _8553_/A _5453_/B _6557_/B _8547_/A vssd1 vssd1 vccd1 vccd1 _7691_/X sky130_fd_sc_hd__o211a_1
XFILLER_32_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6642_ _6999_/A vssd1 vssd1 vccd1 vccd1 _7370_/A sky130_fd_sc_hd__buf_2
XFILLER_32_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6573_ _6579_/A _6579_/B vssd1 vssd1 vccd1 vccd1 _6735_/A sky130_fd_sc_hd__xor2_1
X_8312_ _8368_/A _8312_/B vssd1 vssd1 vccd1 vccd1 _8312_/Y sky130_fd_sc_hd__nor2_1
X_5524_ _5559_/B _5523_/C _5523_/A vssd1 vssd1 vccd1 vccd1 _5533_/B sky130_fd_sc_hd__a21oi_1
X_8243_ _8365_/A _8243_/B vssd1 vssd1 vccd1 vccd1 _8483_/A sky130_fd_sc_hd__nand2_1
X_5455_ _5455_/A _5455_/B vssd1 vssd1 vccd1 vccd1 _5477_/B sky130_fd_sc_hd__nor2_2
X_4406_ _4406_/A vssd1 vssd1 vccd1 vccd1 _4406_/Y sky130_fd_sc_hd__inv_2
X_8174_ _8172_/Y _8174_/B vssd1 vssd1 vccd1 vccd1 _8258_/B sky130_fd_sc_hd__and2b_1
X_7125_ _7125_/A _7125_/B _7125_/C _7125_/D vssd1 vssd1 vccd1 vccd1 _7154_/C sky130_fd_sc_hd__or4_1
X_5386_ _5426_/A _5432_/A _5389_/A _5386_/D vssd1 vssd1 vccd1 vccd1 _5386_/X sky130_fd_sc_hd__and4bb_1
XFILLER_86_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4337_ _4338_/A vssd1 vssd1 vccd1 vccd1 _4337_/Y sky130_fd_sc_hd__inv_2
X_7056_ _7280_/B _7443_/A _7145_/B _7055_/X vssd1 vssd1 vccd1 vccd1 _7057_/B sky130_fd_sc_hd__a31oi_2
XFILLER_59_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6007_ _6200_/A _6007_/B vssd1 vssd1 vccd1 vccd1 _6188_/B sky130_fd_sc_hd__xnor2_1
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7958_ _7958_/A _8026_/B _7958_/C vssd1 vssd1 vccd1 vccd1 _8025_/A sky130_fd_sc_hd__nand3_1
XFILLER_15_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6909_ _7409_/A _7102_/B vssd1 vssd1 vccd1 vccd1 _6911_/A sky130_fd_sc_hd__nor2_1
X_7889_ _7970_/A _8410_/A vssd1 vssd1 vccd1 vccd1 _7891_/C sky130_fd_sc_hd__xnor2_1
XFILLER_23_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5240_ _5244_/A _5240_/B _5245_/D _5240_/D vssd1 vssd1 vccd1 vccd1 _5240_/X sky130_fd_sc_hd__or4_1
XFILLER_102_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5171_ _5171_/A _5171_/B _5171_/C vssd1 vssd1 vccd1 vccd1 _5175_/D sky130_fd_sc_hd__or3_1
XFILLER_68_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8930_ _8930_/A _4451_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[29] sky130_fd_sc_hd__ebufn_8
X_8861_ _8861_/A _4369_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[30] sky130_fd_sc_hd__ebufn_8
XFILLER_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7812_ _7923_/A _7923_/B vssd1 vssd1 vccd1 vccd1 _7819_/A sky130_fd_sc_hd__xor2_1
X_4955_ _4955_/A vssd1 vssd1 vccd1 vccd1 _5091_/C sky130_fd_sc_hd__clkbuf_2
X_7743_ _7905_/B vssd1 vssd1 vccd1 vccd1 _8304_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4886_ _5121_/A _5222_/B vssd1 vssd1 vccd1 vccd1 _4964_/B sky130_fd_sc_hd__or2_1
X_7674_ _8281_/B _7661_/C _8281_/A vssd1 vssd1 vccd1 vccd1 _7675_/B sky130_fd_sc_hd__a21oi_1
X_6625_ _6656_/B vssd1 vssd1 vccd1 vccd1 _6625_/X sky130_fd_sc_hd__clkbuf_2
X_6556_ _6745_/A vssd1 vssd1 vccd1 vccd1 _6558_/A sky130_fd_sc_hd__inv_2
X_5507_ _5521_/B vssd1 vssd1 vccd1 vccd1 _5993_/A sky130_fd_sc_hd__clkbuf_2
X_6487_ _6531_/A vssd1 vssd1 vccd1 vccd1 _6498_/A sky130_fd_sc_hd__inv_2
X_8226_ _8126_/A _8224_/Y _8415_/A vssd1 vssd1 vccd1 vccd1 _8328_/A sky130_fd_sc_hd__o21a_1
X_5438_ _8605_/Q _8668_/Q vssd1 vssd1 vccd1 vccd1 _5439_/A sky130_fd_sc_hd__or2b_1
X_8157_ _8158_/A _8158_/B vssd1 vssd1 vccd1 vccd1 _8256_/A sky130_fd_sc_hd__and2_1
X_5369_ _8669_/Q vssd1 vssd1 vccd1 vccd1 _6341_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7108_ _7125_/B _7125_/C _7125_/D _7107_/X vssd1 vssd1 vccd1 vccd1 _7113_/A sky130_fd_sc_hd__o31a_1
X_8088_ _8087_/A _8087_/B _8087_/C vssd1 vssd1 vccd1 vccd1 _8089_/B sky130_fd_sc_hd__a21oi_1
X_7039_ _7039_/A _7303_/A vssd1 vssd1 vccd1 vccd1 _7040_/B sky130_fd_sc_hd__xor2_1
XFILLER_87_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4740_ _7614_/A _4740_/B vssd1 vssd1 vccd1 vccd1 _4740_/X sky130_fd_sc_hd__or2_1
X_4671_ _4723_/B vssd1 vssd1 vccd1 vccd1 _4727_/A sky130_fd_sc_hd__clkbuf_2
X_6410_ _6413_/B _6410_/B _6464_/B vssd1 vssd1 vccd1 vccd1 _6411_/A sky130_fd_sc_hd__and3b_1
X_7390_ _7390_/A _7390_/B vssd1 vssd1 vccd1 vccd1 _7391_/B sky130_fd_sc_hd__xnor2_1
X_6341_ _6341_/A _8655_/Q vssd1 vssd1 vccd1 vccd1 _6342_/B sky130_fd_sc_hd__or2b_1
XFILLER_103_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6272_ _5746_/B _5974_/B _6195_/B _5952_/B vssd1 vssd1 vccd1 vccd1 _6274_/A sky130_fd_sc_hd__a211o_1
X_5223_ _5223_/A _5223_/B _5230_/B _5223_/D vssd1 vssd1 vccd1 vccd1 _5224_/C sky130_fd_sc_hd__or4_1
X_8011_ _8021_/A _8011_/B _8011_/C vssd1 vssd1 vccd1 vccd1 _8021_/B sky130_fd_sc_hd__nand3_1
XFILLER_102_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5154_ _5154_/A _5154_/B _5154_/C _5224_/B vssd1 vssd1 vccd1 vccd1 _5154_/X sky130_fd_sc_hd__or4_1
XFILLER_69_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5085_ _5175_/A _5091_/C _5208_/A _5244_/C _5084_/X vssd1 vssd1 vccd1 vccd1 _5085_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_56_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8913_ _8913_/A _4428_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[12] sky130_fd_sc_hd__ebufn_8
XFILLER_2_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8844_ _8844_/A _4349_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[13] sky130_fd_sc_hd__ebufn_8
XFILLER_25_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5987_ _5987_/A _5987_/B vssd1 vssd1 vccd1 vccd1 _6191_/B sky130_fd_sc_hd__xnor2_1
X_4938_ _5222_/A _5100_/A vssd1 vssd1 vccd1 vccd1 _5192_/D sky130_fd_sc_hd__nand2_1
X_7726_ _8054_/A _7670_/S _7724_/Y _7725_/Y _7672_/X vssd1 vssd1 vccd1 vccd1 _7727_/B
+ sky130_fd_sc_hd__a32o_1
X_4869_ _4786_/C _4864_/X _4960_/B _4868_/Y vssd1 vssd1 vccd1 vccd1 _5190_/B sky130_fd_sc_hd__a211o_1
X_7657_ _7661_/A vssd1 vssd1 vccd1 vccd1 _7813_/A sky130_fd_sc_hd__clkbuf_2
X_6608_ _6730_/A _6730_/B _7332_/A vssd1 vssd1 vccd1 vccd1 _6617_/A sky130_fd_sc_hd__a21oi_2
XFILLER_21_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7588_ _7630_/A _7584_/X _7587_/Y vssd1 vssd1 vccd1 vccd1 _8718_/D sky130_fd_sc_hd__o21a_1
X_6539_ _6533_/Y _5308_/X _6508_/A _6538_/X vssd1 vssd1 vccd1 vccd1 _8703_/D sky130_fd_sc_hd__a22oi_1
X_8209_ _8450_/B _8442_/A _8388_/A vssd1 vssd1 vccd1 vccd1 _8211_/C sky130_fd_sc_hd__o21a_1
XFILLER_101_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5910_ _6030_/A _5910_/B vssd1 vssd1 vccd1 vccd1 _6242_/A sky130_fd_sc_hd__nand2_2
X_6890_ _6890_/A _7350_/A vssd1 vssd1 vccd1 vccd1 _6958_/A sky130_fd_sc_hd__or2_1
XFILLER_19_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5841_ _5841_/A vssd1 vssd1 vccd1 vccd1 _5842_/A sky130_fd_sc_hd__inv_2
XFILLER_61_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8560_ _8576_/A _8560_/B vssd1 vssd1 vccd1 vccd1 _8561_/B sky130_fd_sc_hd__and2b_1
X_5772_ _5727_/A _5772_/B vssd1 vssd1 vccd1 vccd1 _5772_/X sky130_fd_sc_hd__and2b_1
XFILLER_34_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4723_ _4726_/B _4723_/B _4723_/C vssd1 vssd1 vccd1 vccd1 _4724_/A sky130_fd_sc_hd__and3b_1
X_7511_ _7499_/X _8708_/Q _7497_/X _7510_/X vssd1 vssd1 vccd1 vccd1 _8708_/D sky130_fd_sc_hd__o22a_1
X_8491_ _8491_/A _8491_/B vssd1 vssd1 vccd1 vccd1 _8492_/B sky130_fd_sc_hd__xnor2_1
X_7442_ _7372_/A _7372_/B _7376_/A vssd1 vssd1 vccd1 vccd1 _7445_/A sky130_fd_sc_hd__a21bo_1
X_4654_ _5222_/A vssd1 vssd1 vccd1 vccd1 _4923_/A sky130_fd_sc_hd__clkbuf_2
X_7373_ _7447_/D _7373_/B _7373_/C vssd1 vssd1 vccd1 vccd1 _7376_/A sky130_fd_sc_hd__nand3_1
X_4585_ _4607_/A vssd1 vssd1 vccd1 vccd1 _4612_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6324_ _6336_/A _6320_/X _6323_/X _7537_/B vssd1 vssd1 vccd1 vccd1 _6324_/X sky130_fd_sc_hd__o31a_1
X_6255_ _6255_/A _6255_/B vssd1 vssd1 vccd1 vccd1 _6258_/A sky130_fd_sc_hd__or2_1
X_5206_ _5065_/A _5171_/C _5198_/X _5205_/X _5080_/Y vssd1 vssd1 vccd1 vccd1 _5206_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_57_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6186_ _6186_/A _6186_/B vssd1 vssd1 vccd1 vccd1 _6231_/A sky130_fd_sc_hd__xnor2_4
X_5137_ _5223_/D _5230_/D _5231_/D vssd1 vssd1 vccd1 vccd1 _5137_/X sky130_fd_sc_hd__o21a_1
XFILLER_96_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5068_ _5193_/B _5096_/C _5067_/Y vssd1 vssd1 vccd1 vccd1 _5068_/Y sky130_fd_sc_hd__nor3b_1
XFILLER_16_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8771__38 vssd1 vssd1 vccd1 vccd1 _8771__38/HI _8866_/A sky130_fd_sc_hd__conb_1
XFILLER_40_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7709_ _8122_/C vssd1 vssd1 vccd1 vccd1 _8124_/A sky130_fd_sc_hd__buf_2
X_8689_ _8689_/CLK _8689_/D vssd1 vssd1 vccd1 vccd1 _8689_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4370_ _4370_/A vssd1 vssd1 vccd1 vccd1 _4375_/A sky130_fd_sc_hd__buf_6
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6040_ _6063_/A _6063_/B vssd1 vssd1 vccd1 vccd1 _6040_/Y sky130_fd_sc_hd__nand2_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7991_ _8167_/A _8378_/A vssd1 vssd1 vccd1 vccd1 _7998_/A sky130_fd_sc_hd__xor2_2
X_6942_ _6949_/A _6949_/B vssd1 vssd1 vccd1 vccd1 _6944_/B sky130_fd_sc_hd__xor2_1
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6873_ _7371_/A vssd1 vssd1 vccd1 vccd1 _7355_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_62_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8612_ _8671_/CLK _8612_/D vssd1 vssd1 vccd1 vccd1 _8612_/Q sky130_fd_sc_hd__dfxtp_1
X_5824_ _5824_/A _5824_/B vssd1 vssd1 vccd1 vccd1 _5825_/B sky130_fd_sc_hd__nor2_1
XFILLER_22_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5755_ _5845_/A _5755_/B vssd1 vssd1 vccd1 vccd1 _5756_/B sky130_fd_sc_hd__nor2_1
X_8543_ _8542_/Y _8540_/A _8543_/S vssd1 vssd1 vccd1 vccd1 _8544_/B sky130_fd_sc_hd__mux2_1
X_4706_ _5229_/A vssd1 vssd1 vccd1 vccd1 _5053_/A sky130_fd_sc_hd__clkbuf_2
X_8474_ _8474_/A _8474_/B vssd1 vssd1 vccd1 vccd1 _8476_/A sky130_fd_sc_hd__or2_1
X_5686_ _6049_/B _5686_/B vssd1 vssd1 vccd1 vccd1 _5687_/B sky130_fd_sc_hd__nor2_1
X_7425_ _7425_/A _7425_/B vssd1 vssd1 vccd1 vccd1 _7428_/A sky130_fd_sc_hd__xnor2_1
X_4637_ _8598_/Q _8597_/Q _4637_/C vssd1 vssd1 vccd1 vccd1 _4643_/C sky130_fd_sc_hd__and3_1
X_7356_ _7356_/A vssd1 vssd1 vccd1 vccd1 _7455_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4568_ _4568_/A vssd1 vssd1 vccd1 vccd1 _8883_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_103_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7287_ _7266_/X _7473_/B _7472_/A vssd1 vssd1 vccd1 vccd1 _7481_/B sky130_fd_sc_hd__a21oi_2
X_6307_ _6307_/A _6307_/B vssd1 vssd1 vccd1 vccd1 _6309_/A sky130_fd_sc_hd__xnor2_1
X_4499_ _8617_/Q vssd1 vssd1 vccd1 vccd1 _5591_/A sky130_fd_sc_hd__buf_2
X_6238_ _6238_/A _6238_/B vssd1 vssd1 vccd1 vccd1 _6282_/A sky130_fd_sc_hd__xnor2_2
XFILLER_76_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8816__83 vssd1 vssd1 vccd1 vccd1 _8816__83/HI _8925_/A sky130_fd_sc_hd__conb_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6169_ _5955_/A _5955_/B _6168_/X vssd1 vssd1 vccd1 vccd1 _6178_/A sky130_fd_sc_hd__a21bo_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5540_ _5540_/A _6316_/A vssd1 vssd1 vccd1 vccd1 _5560_/A sky130_fd_sc_hd__xnor2_2
X_5471_ _5493_/A _5471_/B vssd1 vssd1 vccd1 vccd1 _5519_/A sky130_fd_sc_hd__nand2_1
X_7210_ _7210_/A _7210_/B vssd1 vssd1 vccd1 vccd1 _7233_/A sky130_fd_sc_hd__xnor2_1
X_4422_ _4425_/A vssd1 vssd1 vccd1 vccd1 _4422_/Y sky130_fd_sc_hd__inv_2
X_8190_ _8190_/A _8164_/B vssd1 vssd1 vccd1 vccd1 _8190_/X sky130_fd_sc_hd__or2b_1
X_4353_ _4357_/A vssd1 vssd1 vccd1 vccd1 _4353_/Y sky130_fd_sc_hd__inv_2
X_7141_ _7141_/A _7141_/B _7141_/C vssd1 vssd1 vccd1 vccd1 _7143_/B sky130_fd_sc_hd__nand3_1
X_7072_ _7072_/A _7072_/B vssd1 vssd1 vccd1 vccd1 _7072_/X sky130_fd_sc_hd__or2_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6023_ _5872_/B _5575_/A _5556_/A _5554_/X vssd1 vssd1 vccd1 vccd1 _6024_/C sky130_fd_sc_hd__a22o_1
XFILLER_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7974_ _8045_/A _8045_/B vssd1 vssd1 vccd1 vccd1 _7975_/B sky130_fd_sc_hd__xor2_1
X_6925_ _6818_/A _6818_/B _6924_/Y vssd1 vssd1 vccd1 vccd1 _6940_/A sky130_fd_sc_hd__a21o_1
XFILLER_22_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6856_ _6856_/A _6856_/B vssd1 vssd1 vccd1 vccd1 _6859_/A sky130_fd_sc_hd__xnor2_1
XFILLER_50_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6787_ _6869_/A _6869_/B vssd1 vssd1 vccd1 vccd1 _6789_/C sky130_fd_sc_hd__xnor2_1
XFILLER_10_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5807_ _5868_/A _5807_/B vssd1 vssd1 vccd1 vccd1 _5808_/B sky130_fd_sc_hd__and2_1
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5738_ _5738_/A _6238_/A vssd1 vssd1 vccd1 vccd1 _5751_/C sky130_fd_sc_hd__xnor2_1
XFILLER_22_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8526_ _8531_/A _8726_/Q vssd1 vssd1 vccd1 vccd1 _8526_/Y sky130_fd_sc_hd__nor2_1
X_5669_ _5669_/A _5669_/B vssd1 vssd1 vccd1 vccd1 _5691_/B sky130_fd_sc_hd__nand2_1
X_8457_ _8411_/S _8412_/A _8456_/X vssd1 vssd1 vccd1 vccd1 _8459_/A sky130_fd_sc_hd__a21bo_1
X_7408_ _7316_/A _7316_/B _7315_/A vssd1 vssd1 vccd1 vccd1 _7412_/A sky130_fd_sc_hd__o21ai_1
XFILLER_2_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8388_ _8388_/A _8327_/B vssd1 vssd1 vccd1 vccd1 _8392_/B sky130_fd_sc_hd__or2b_1
X_7339_ _7339_/A _7339_/B vssd1 vssd1 vccd1 vccd1 _7419_/B sky130_fd_sc_hd__xnor2_1
XFILLER_89_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_2_1_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_95_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4971_ _4946_/X _4959_/X _4960_/X _4970_/X vssd1 vssd1 vccd1 vccd1 _4971_/X sky130_fd_sc_hd__o31a_1
XFILLER_63_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6710_ _6710_/A _6774_/S vssd1 vssd1 vccd1 vccd1 _7369_/A sky130_fd_sc_hd__xnor2_2
XFILLER_51_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7690_ _8731_/Q vssd1 vssd1 vccd1 vccd1 _8547_/A sky130_fd_sc_hd__inv_2
X_6641_ _7000_/A vssd1 vssd1 vccd1 vccd1 _6999_/A sky130_fd_sc_hd__buf_2
X_6572_ _8700_/Q _8617_/Q vssd1 vssd1 vccd1 vccd1 _6579_/B sky130_fd_sc_hd__xnor2_4
X_8311_ _8311_/A _8370_/B vssd1 vssd1 vccd1 vccd1 _8489_/B sky130_fd_sc_hd__xnor2_2
X_5523_ _5523_/A _5559_/B _5523_/C vssd1 vssd1 vccd1 vccd1 _5533_/A sky130_fd_sc_hd__and3_1
X_8242_ _8378_/A _8242_/B vssd1 vssd1 vccd1 vccd1 _8278_/A sky130_fd_sc_hd__nand2_1
X_5454_ _5453_/B _8671_/Q vssd1 vssd1 vccd1 vccd1 _5455_/B sky130_fd_sc_hd__and2b_1
X_4405_ _4406_/A vssd1 vssd1 vccd1 vccd1 _4405_/Y sky130_fd_sc_hd__inv_2
X_8173_ _8172_/A _8172_/C _8172_/B vssd1 vssd1 vccd1 vccd1 _8174_/B sky130_fd_sc_hd__o21ai_1
X_5385_ _5404_/B _5400_/A _5411_/B vssd1 vssd1 vccd1 vccd1 _5386_/D sky130_fd_sc_hd__o21ai_1
X_7124_ _7107_/A _7127_/B _7124_/C _7124_/D vssd1 vssd1 vccd1 vccd1 _7125_/A sky130_fd_sc_hd__and4bb_1
X_4336_ _4338_/A vssd1 vssd1 vccd1 vccd1 _4336_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7055_ _7335_/A _7196_/C _6797_/A vssd1 vssd1 vccd1 vccd1 _7055_/X sky130_fd_sc_hd__o21a_1
XFILLER_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6006_ _6006_/A _6199_/A vssd1 vssd1 vccd1 vccd1 _6007_/B sky130_fd_sc_hd__xnor2_1
XFILLER_67_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7957_ _7956_/B _8026_/A _8123_/S vssd1 vssd1 vccd1 vccd1 _7958_/C sky130_fd_sc_hd__a21bo_1
X_6908_ _6802_/A _6802_/B _6907_/X vssd1 vssd1 vccd1 vccd1 _6995_/A sky130_fd_sc_hd__a21oi_1
X_7888_ _7888_/A vssd1 vssd1 vccd1 vccd1 _8410_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_42_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6839_ _7060_/A _6839_/B vssd1 vssd1 vccd1 vccd1 _7145_/A sky130_fd_sc_hd__nor2_2
XFILLER_50_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8509_ _8509_/A _8509_/B _8509_/C vssd1 vssd1 vccd1 vccd1 _8510_/B sky130_fd_sc_hd__and3_1
XFILLER_2_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5170_ _5208_/A _5170_/B vssd1 vssd1 vccd1 vccd1 _5240_/D sky130_fd_sc_hd__or2_1
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8860_ _8860_/A _4368_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[29] sky130_fd_sc_hd__ebufn_8
XFILLER_64_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7811_ _8281_/A _7661_/X _7748_/Y _7662_/A vssd1 vssd1 vccd1 vccd1 _7923_/B sky130_fd_sc_hd__a211o_1
XFILLER_36_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4954_ _4916_/A _5222_/D _4941_/X _4953_/X vssd1 vssd1 vccd1 vccd1 _4954_/X sky130_fd_sc_hd__o31a_1
XFILLER_51_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7742_ _7742_/A _7742_/B vssd1 vssd1 vccd1 vccd1 _7905_/B sky130_fd_sc_hd__xnor2_2
X_4885_ _4891_/A _4885_/B _4891_/C vssd1 vssd1 vccd1 vccd1 _5222_/B sky130_fd_sc_hd__nor3_1
XFILLER_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7673_ _7736_/A _7671_/B _7672_/X vssd1 vssd1 vccd1 vccd1 _7675_/A sky130_fd_sc_hd__a21bo_1
X_6624_ _6639_/A _8621_/Q vssd1 vssd1 vccd1 vccd1 _6656_/B sky130_fd_sc_hd__or2_1
X_6555_ _6557_/B _8711_/Q vssd1 vssd1 vccd1 vccd1 _6745_/A sky130_fd_sc_hd__or2b_1
X_5506_ _5506_/A _5506_/B vssd1 vssd1 vccd1 vccd1 _5521_/B sky130_fd_sc_hd__and2_1
X_6486_ _8702_/Q vssd1 vssd1 vccd1 vccd1 _6531_/A sky130_fd_sc_hd__clkbuf_2
X_8225_ _8225_/A vssd1 vssd1 vccd1 vccd1 _8415_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5437_ _5437_/A vssd1 vssd1 vccd1 vccd1 _8663_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8156_ _8200_/A _8156_/B vssd1 vssd1 vccd1 vccd1 _8158_/B sky130_fd_sc_hd__and2_1
X_5368_ _8670_/Q vssd1 vssd1 vccd1 vccd1 _5456_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5299_ _5299_/A vssd1 vssd1 vccd1 vccd1 _8634_/D sky130_fd_sc_hd__clkbuf_1
X_7107_ _7107_/A _7127_/B _7124_/C _7124_/D vssd1 vssd1 vccd1 vccd1 _7107_/X sky130_fd_sc_hd__or4bb_1
XFILLER_59_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8087_ _8087_/A _8087_/B _8087_/C vssd1 vssd1 vccd1 vccd1 _8258_/A sky130_fd_sc_hd__and3_1
XFILLER_101_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7038_ _7304_/A _7304_/B vssd1 vssd1 vccd1 vccd1 _7303_/A sky130_fd_sc_hd__xnor2_1
XFILLER_101_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8777__44 vssd1 vssd1 vccd1 vccd1 _8777__44/HI _8872_/A sky130_fd_sc_hd__conb_1
XFILLER_46_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4670_ _5296_/A _4752_/A vssd1 vssd1 vccd1 vccd1 _4723_/B sky130_fd_sc_hd__and2_1
X_6340_ _8655_/Q _6341_/A vssd1 vssd1 vccd1 vccd1 _6342_/A sky130_fd_sc_hd__or2b_1
XFILLER_6_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6271_ _6176_/A _6176_/B _6270_/X vssd1 vssd1 vccd1 vccd1 _6275_/A sky130_fd_sc_hd__a21oi_1
X_5222_ _5222_/A _5222_/B _5223_/B _5222_/D vssd1 vssd1 vccd1 vccd1 _5222_/X sky130_fd_sc_hd__or4_1
X_8010_ _8020_/A _8020_/B vssd1 vssd1 vccd1 vccd1 _8011_/C sky130_fd_sc_hd__xor2_1
X_5153_ _5153_/A _5153_/B vssd1 vssd1 vccd1 vccd1 _5153_/X sky130_fd_sc_hd__and2_1
XFILLER_69_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5084_ _5199_/A _5207_/B _5084_/C vssd1 vssd1 vccd1 vccd1 _5084_/X sky130_fd_sc_hd__or3_1
X_8912_ _8912_/A _4425_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[11] sky130_fd_sc_hd__ebufn_8
XFILLER_71_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8843_ _8843_/A _4348_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[12] sky130_fd_sc_hd__ebufn_8
XFILLER_37_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5986_ _6211_/B _5986_/B vssd1 vssd1 vccd1 vccd1 _5987_/B sky130_fd_sc_hd__xnor2_1
X_4937_ _4937_/A _4937_/B vssd1 vssd1 vccd1 vccd1 _5100_/A sky130_fd_sc_hd__or2_1
X_7725_ _7725_/A _7725_/B vssd1 vssd1 vccd1 vccd1 _7725_/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7656_ _7656_/A _7656_/B vssd1 vssd1 vccd1 vccd1 _7661_/A sky130_fd_sc_hd__xor2_2
X_4868_ _4868_/A _4896_/A vssd1 vssd1 vccd1 vccd1 _4868_/Y sky130_fd_sc_hd__nor2_1
X_6607_ _6607_/A vssd1 vssd1 vccd1 vccd1 _7332_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4799_ _4799_/A _4859_/A _4899_/B _4799_/D vssd1 vssd1 vccd1 vccd1 _4799_/X sky130_fd_sc_hd__or4_1
X_7587_ _7630_/A _8574_/A _7544_/X vssd1 vssd1 vccd1 vccd1 _7587_/Y sky130_fd_sc_hd__a21oi_1
X_6538_ _6538_/A _6538_/B vssd1 vssd1 vccd1 vccd1 _6538_/X sky130_fd_sc_hd__xor2_1
X_6469_ _8651_/Q _8650_/Q vssd1 vssd1 vccd1 vccd1 _6471_/C sky130_fd_sc_hd__nor2_1
X_8208_ _8208_/A _8450_/B vssd1 vssd1 vccd1 vccd1 _8388_/A sky130_fd_sc_hd__nand2_2
X_8139_ _8139_/A _8139_/B vssd1 vssd1 vccd1 vccd1 _8450_/B sky130_fd_sc_hd__nor2_2
XFILLER_101_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5840_ _5838_/Y _5840_/B vssd1 vssd1 vccd1 vccd1 _5924_/B sky130_fd_sc_hd__and2b_1
XFILLER_34_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5771_ _6018_/A _6018_/B _5770_/X vssd1 vssd1 vccd1 vccd1 _5851_/A sky130_fd_sc_hd__a21o_1
X_4722_ _4711_/A _4715_/A _6746_/B vssd1 vssd1 vccd1 vccd1 _4723_/C sky130_fd_sc_hd__o21ai_1
X_7510_ _7510_/A _7510_/B _7510_/C vssd1 vssd1 vccd1 vccd1 _7510_/X sky130_fd_sc_hd__and3_1
X_8490_ _8490_/A _8490_/B vssd1 vssd1 vccd1 vccd1 _8491_/B sky130_fd_sc_hd__xnor2_1
X_7441_ _7441_/A _7441_/B vssd1 vssd1 vccd1 vccd1 _7458_/A sky130_fd_sc_hd__xnor2_1
X_4653_ _5245_/A vssd1 vssd1 vccd1 vccd1 _5222_/A sky130_fd_sc_hd__clkbuf_2
X_7372_ _7372_/A _7372_/B vssd1 vssd1 vccd1 vccd1 _7373_/C sky130_fd_sc_hd__xor2_1
X_4584_ _6503_/A _8601_/Q vssd1 vssd1 vccd1 vccd1 _4607_/A sky130_fd_sc_hd__nor2_1
X_6323_ _6297_/A _6332_/C _6300_/X _6296_/X vssd1 vssd1 vccd1 vccd1 _6323_/X sky130_fd_sc_hd__a211o_1
X_6254_ _6209_/A _6207_/X _6253_/X vssd1 vssd1 vccd1 vccd1 _6259_/A sky130_fd_sc_hd__o21a_1
XFILLER_103_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5205_ _5205_/A _5205_/B _5205_/C vssd1 vssd1 vccd1 vccd1 _5205_/X sky130_fd_sc_hd__or3_1
X_6185_ _6185_/A vssd1 vssd1 vccd1 vccd1 _6186_/B sky130_fd_sc_hd__clkinv_2
XFILLER_96_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5136_ _5245_/A _5136_/B _5136_/C vssd1 vssd1 vccd1 vccd1 _5231_/D sky130_fd_sc_hd__or3_1
XFILLER_57_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5067_ _5175_/B _5084_/C _5067_/C vssd1 vssd1 vccd1 vccd1 _5067_/Y sky130_fd_sc_hd__nor3_1
XFILLER_84_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5969_ _6172_/A _5969_/B vssd1 vssd1 vccd1 vccd1 _5976_/A sky130_fd_sc_hd__xnor2_2
XFILLER_12_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7708_ _7955_/A vssd1 vssd1 vccd1 vccd1 _8122_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_8688_ _8689_/CLK _8688_/D vssd1 vssd1 vccd1 vccd1 _8688_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7639_ _7639_/A _7639_/B vssd1 vssd1 vccd1 vccd1 _7834_/A sky130_fd_sc_hd__xnor2_2
XFILLER_4_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8747__14 vssd1 vssd1 vccd1 vccd1 _8747__14/HI _8842_/A sky130_fd_sc_hd__conb_1
XFILLER_56_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7990_ _7990_/A vssd1 vssd1 vccd1 vccd1 _8378_/A sky130_fd_sc_hd__buf_2
XFILLER_26_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6941_ _6941_/A _7047_/A vssd1 vssd1 vccd1 vccd1 _6949_/B sky130_fd_sc_hd__xor2_1
XFILLER_81_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6872_ _6872_/A _6892_/A vssd1 vssd1 vccd1 vccd1 _7371_/A sky130_fd_sc_hd__xnor2_1
XFILLER_81_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8611_ _8671_/CLK _8611_/D vssd1 vssd1 vccd1 vccd1 _8611_/Q sky130_fd_sc_hd__dfxtp_1
X_5823_ _5824_/A _5824_/B vssd1 vssd1 vccd1 vccd1 _5922_/A sky130_fd_sc_hd__and2_1
XFILLER_22_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8542_ _8729_/Q _8542_/B vssd1 vssd1 vccd1 vccd1 _8542_/Y sky130_fd_sc_hd__xnor2_1
X_5754_ _5754_/A _5754_/B _5754_/C vssd1 vssd1 vccd1 vccd1 _5755_/B sky130_fd_sc_hd__and3_1
X_4705_ _8604_/Q vssd1 vssd1 vccd1 vccd1 _5229_/A sky130_fd_sc_hd__inv_2
X_8473_ _8312_/B _8310_/B _8473_/S vssd1 vssd1 vccd1 vccd1 _8474_/B sky130_fd_sc_hd__mux2_1
X_5685_ _5685_/A _5685_/B vssd1 vssd1 vccd1 vccd1 _5686_/B sky130_fd_sc_hd__and2_1
X_7424_ _7424_/A _7424_/B vssd1 vssd1 vccd1 vccd1 _7425_/B sky130_fd_sc_hd__xnor2_1
X_4636_ _8597_/Q _4637_/C _4635_/Y vssd1 vssd1 vccd1 vccd1 _8597_/D sky130_fd_sc_hd__a21oi_1
X_7355_ _7355_/A _7355_/B _7355_/C vssd1 vssd1 vccd1 vccd1 _7356_/A sky130_fd_sc_hd__or3_1
X_4567_ _8629_/Q _4567_/B vssd1 vssd1 vccd1 vccd1 _4568_/A sky130_fd_sc_hd__and2_1
X_6306_ _6306_/A _6306_/B vssd1 vssd1 vccd1 vccd1 _6306_/X sky130_fd_sc_hd__xor2_1
XFILLER_89_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4498_ _4864_/A vssd1 vssd1 vccd1 vccd1 _4799_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7286_ _7286_/A _7286_/B _7286_/C vssd1 vssd1 vccd1 vccd1 _7472_/A sky130_fd_sc_hd__and3_1
XFILLER_89_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6237_ _6302_/A _6302_/B _6312_/B _6236_/Y _6235_/B vssd1 vssd1 vccd1 vccd1 _6294_/A
+ sky130_fd_sc_hd__a32o_2
XFILLER_85_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6168_ _6168_/A _5954_/B vssd1 vssd1 vccd1 vccd1 _6168_/X sky130_fd_sc_hd__or2b_1
XFILLER_94_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5119_ _5119_/A _5245_/C vssd1 vssd1 vccd1 vccd1 _5227_/C sky130_fd_sc_hd__or2_2
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6099_ _6119_/A _6119_/B _6099_/C vssd1 vssd1 vccd1 vccd1 _6101_/A sky130_fd_sc_hd__and3_1
XFILLER_27_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_3_3_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_7_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_25_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5470_ _5470_/A _6598_/A vssd1 vssd1 vccd1 vccd1 _5471_/B sky130_fd_sc_hd__nand2_1
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4421_ _4425_/A vssd1 vssd1 vccd1 vccd1 _4421_/Y sky130_fd_sc_hd__inv_2
X_4352_ _4370_/A vssd1 vssd1 vccd1 vccd1 _4357_/A sky130_fd_sc_hd__clkbuf_2
X_7140_ _7181_/A _7181_/B _7139_/C vssd1 vssd1 vccd1 vccd1 _7141_/C sky130_fd_sc_hd__a21o_1
X_7071_ _7147_/B _7167_/A _7147_/A vssd1 vssd1 vccd1 vccd1 _7148_/A sky130_fd_sc_hd__o21a_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6022_ _6069_/A _6069_/B vssd1 vssd1 vccd1 vccd1 _6024_/B sky130_fd_sc_hd__and2b_1
XFILLER_39_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7973_ _8044_/A _7973_/B vssd1 vssd1 vccd1 vccd1 _8045_/B sky130_fd_sc_hd__xnor2_1
X_6924_ _6924_/A _6924_/B vssd1 vssd1 vccd1 vccd1 _6924_/Y sky130_fd_sc_hd__nor2_1
XFILLER_81_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6855_ _6926_/A _6926_/B vssd1 vssd1 vccd1 vccd1 _6856_/B sky130_fd_sc_hd__xnor2_2
X_6786_ _6905_/A _6786_/B vssd1 vssd1 vccd1 vccd1 _6869_/B sky130_fd_sc_hd__xnor2_2
XFILLER_50_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5806_ _5806_/A _5806_/B _6209_/A vssd1 vssd1 vccd1 vccd1 _5807_/B sky130_fd_sc_hd__nand3_1
X_5737_ _5737_/A _5816_/A vssd1 vssd1 vccd1 vccd1 _6238_/A sky130_fd_sc_hd__xnor2_4
XFILLER_22_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8525_ _8525_/A _8525_/B _8529_/B _8525_/D vssd1 vssd1 vccd1 vccd1 _8525_/X sky130_fd_sc_hd__or4_1
X_8456_ _8399_/A _8139_/B _8411_/S _8412_/A _8412_/B vssd1 vssd1 vccd1 vccd1 _8456_/X
+ sky130_fd_sc_hd__a32o_1
X_7407_ _7322_/A _7322_/B _7406_/X vssd1 vssd1 vccd1 vccd1 _7424_/A sky130_fd_sc_hd__a21oi_1
XFILLER_89_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5668_ _5669_/A _5669_/B vssd1 vssd1 vccd1 vccd1 _5754_/B sky130_fd_sc_hd__or2_1
X_4619_ _8592_/Q _8591_/Q _4619_/C vssd1 vssd1 vccd1 vccd1 _4623_/B sky130_fd_sc_hd__and3_1
X_8387_ _8387_/A _8326_/A vssd1 vssd1 vccd1 vccd1 _8392_/A sky130_fd_sc_hd__or2b_1
X_5599_ _8660_/Q _7643_/B vssd1 vssd1 vccd1 vccd1 _5599_/X sky130_fd_sc_hd__and2b_1
XFILLER_104_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7338_ _7338_/A _7338_/B vssd1 vssd1 vccd1 vccd1 _7339_/B sky130_fd_sc_hd__xor2_2
XFILLER_2_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7269_ _7269_/A vssd1 vssd1 vccd1 vccd1 _7272_/B sky130_fd_sc_hd__inv_2
XFILLER_77_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4970_ _5190_/B _4970_/B _4970_/C _5139_/C vssd1 vssd1 vccd1 vccd1 _4970_/X sky130_fd_sc_hd__or4_1
XFILLER_17_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6640_ _6625_/X _6688_/A _6689_/A _6690_/A _7082_/A vssd1 vssd1 vccd1 vccd1 _7000_/A
+ sky130_fd_sc_hd__a311o_4
XFILLER_32_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6571_ _6588_/A _6578_/B _6570_/X vssd1 vssd1 vccd1 vccd1 _6579_/A sky130_fd_sc_hd__a21o_1
X_8310_ _8312_/B _8310_/B vssd1 vssd1 vccd1 vccd1 _8370_/B sky130_fd_sc_hd__and2_2
X_5522_ _5874_/A _5521_/B _5521_/C _5559_/A vssd1 vssd1 vccd1 vccd1 _5523_/C sky130_fd_sc_hd__a22o_1
X_8241_ _8274_/A _8274_/B vssd1 vssd1 vccd1 vccd1 _8260_/A sky130_fd_sc_hd__xor2_2
X_5453_ _8671_/Q _5453_/B vssd1 vssd1 vccd1 vccd1 _5455_/A sky130_fd_sc_hd__and2b_1
X_4404_ _4406_/A vssd1 vssd1 vccd1 vccd1 _4404_/Y sky130_fd_sc_hd__inv_2
X_5384_ _8660_/Q vssd1 vssd1 vccd1 vccd1 _5411_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_8172_ _8172_/A _8172_/B _8172_/C vssd1 vssd1 vccd1 vccd1 _8172_/Y sky130_fd_sc_hd__nor3_1
XFILLER_99_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7123_ _7395_/A _7395_/B vssd1 vssd1 vccd1 vccd1 _7488_/A sky130_fd_sc_hd__xor2_2
X_4335_ _4338_/A vssd1 vssd1 vccd1 vccd1 _4335_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7054_ _7430_/A _7054_/B vssd1 vssd1 vccd1 vccd1 _7145_/B sky130_fd_sc_hd__nor2_2
X_6005_ _6005_/A _6005_/B vssd1 vssd1 vccd1 vccd1 _6199_/A sky130_fd_sc_hd__xnor2_1
XFILLER_55_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8801__68 vssd1 vssd1 vccd1 vccd1 _8801__68/HI _8910_/A sky130_fd_sc_hd__conb_1
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7956_ _8123_/S _7956_/B _8026_/A vssd1 vssd1 vccd1 vccd1 _8026_/B sky130_fd_sc_hd__nand3b_1
XFILLER_42_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6907_ _6801_/A _6907_/B vssd1 vssd1 vccd1 vccd1 _6907_/X sky130_fd_sc_hd__and2b_1
X_7887_ _7887_/A _7887_/B vssd1 vssd1 vccd1 vccd1 _7970_/A sky130_fd_sc_hd__nand2_1
XFILLER_35_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6838_ _7009_/B _6927_/A vssd1 vssd1 vccd1 vccd1 _7432_/B sky130_fd_sc_hd__nor2_2
X_6769_ _6769_/A _6728_/B vssd1 vssd1 vccd1 vccd1 _6789_/B sky130_fd_sc_hd__or2b_1
XFILLER_10_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8508_ _8508_/A _8508_/B vssd1 vssd1 vccd1 vccd1 _8508_/Y sky130_fd_sc_hd__nor2_1
X_8439_ _8379_/B _8439_/B vssd1 vssd1 vccd1 vccd1 _8439_/X sky130_fd_sc_hd__and2b_1
XFILLER_2_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7810_ _7901_/A _7901_/B vssd1 vssd1 vccd1 vccd1 _7923_/A sky130_fd_sc_hd__xnor2_1
XFILLER_64_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4953_ _5215_/A _5171_/B _5166_/B _4953_/D vssd1 vssd1 vccd1 vccd1 _4953_/X sky130_fd_sc_hd__or4_1
XFILLER_51_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7741_ _7741_/A _7741_/B vssd1 vssd1 vccd1 vccd1 _7742_/B sky130_fd_sc_hd__nand2_1
XFILLER_51_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7672_ _7725_/A _7725_/B vssd1 vssd1 vccd1 vccd1 _7672_/X sky130_fd_sc_hd__or2_1
X_6623_ _7293_/A vssd1 vssd1 vccd1 vccd1 _7392_/A sky130_fd_sc_hd__clkbuf_2
X_4884_ _4919_/A _4948_/B vssd1 vssd1 vccd1 vccd1 _5121_/A sky130_fd_sc_hd__nor2_1
XFILLER_32_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6554_ _6593_/A _6582_/B _6553_/X vssd1 vssd1 vccd1 vccd1 _6559_/A sky130_fd_sc_hd__a21o_1
XFILLER_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6485_ _6475_/X _6484_/X _8558_/A vssd1 vssd1 vccd1 vccd1 _8696_/D sky130_fd_sc_hd__a21oi_1
X_5505_ _5792_/B vssd1 vssd1 vccd1 vccd1 _5872_/B sky130_fd_sc_hd__clkbuf_2
X_5436_ _7550_/A _5436_/B _5436_/C vssd1 vssd1 vccd1 vccd1 _5437_/A sky130_fd_sc_hd__and3_1
XFILLER_10_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8224_ _8224_/A _8323_/A vssd1 vssd1 vccd1 vccd1 _8224_/Y sky130_fd_sc_hd__nor2_1
X_8155_ _8155_/A _8390_/A vssd1 vssd1 vccd1 vccd1 _8156_/B sky130_fd_sc_hd__or2_1
X_5367_ _5374_/A _5389_/A vssd1 vssd1 vccd1 vccd1 _5367_/Y sky130_fd_sc_hd__nand2_1
XFILLER_101_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5298_ _8634_/Q _5359_/A vssd1 vssd1 vccd1 vccd1 _5299_/A sky130_fd_sc_hd__and2b_1
XFILLER_87_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7106_ _7105_/B _7105_/C _7105_/A vssd1 vssd1 vccd1 vccd1 _7125_/D sky130_fd_sc_hd__a21oi_1
X_8086_ _7813_/A _7998_/A _8308_/A vssd1 vssd1 vccd1 vccd1 _8087_/C sky130_fd_sc_hd__a21oi_1
X_7037_ _6935_/A _6934_/B _6934_/A vssd1 vssd1 vccd1 vccd1 _7304_/B sky130_fd_sc_hd__a21boi_1
XFILLER_74_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7939_ _7940_/A _7940_/B _7940_/C vssd1 vssd1 vccd1 vccd1 _8017_/A sky130_fd_sc_hd__a21oi_1
XFILLER_42_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8792__59 vssd1 vssd1 vccd1 vccd1 _8792__59/HI _8901_/A sky130_fd_sc_hd__conb_1
XFILLER_14_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6270_ _6175_/A _6270_/B vssd1 vssd1 vccd1 vccd1 _6270_/X sky130_fd_sc_hd__and2b_1
XFILLER_102_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5221_ _5179_/B _5218_/X _5220_/X _5080_/A vssd1 vssd1 vccd1 vccd1 _5221_/X sky130_fd_sc_hd__o211a_1
X_5152_ _4795_/B _4702_/A _4661_/A _5150_/X _5151_/X vssd1 vssd1 vccd1 vccd1 _5152_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_69_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5083_ _5096_/A _5056_/Y _5064_/X _5082_/X vssd1 vssd1 vccd1 vccd1 _5083_/X sky130_fd_sc_hd__a31o_1
XFILLER_56_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8911_ _8911_/A _4423_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[10] sky130_fd_sc_hd__ebufn_8
X_8842_ _8842_/A _4347_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[11] sky130_fd_sc_hd__ebufn_8
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7724_ _7835_/A _7813_/A vssd1 vssd1 vccd1 vccd1 _7724_/Y sky130_fd_sc_hd__nand2_1
X_5985_ _5567_/B _5876_/S _5893_/B _5981_/A vssd1 vssd1 vccd1 vccd1 _5986_/B sky130_fd_sc_hd__o2bb2a_1
X_4936_ _4998_/B vssd1 vssd1 vccd1 vccd1 _5245_/B sky130_fd_sc_hd__clkbuf_2
X_4867_ _4899_/B _4867_/B vssd1 vssd1 vccd1 vccd1 _4960_/B sky130_fd_sc_hd__nor2_2
X_7655_ _8515_/A _8145_/A vssd1 vssd1 vccd1 vccd1 _7661_/C sky130_fd_sc_hd__or2_1
X_6606_ _6825_/A _6826_/A _6826_/B _6605_/X vssd1 vssd1 vccd1 vccd1 _6730_/B sky130_fd_sc_hd__a31o_2
X_7586_ _8543_/S vssd1 vssd1 vccd1 vccd1 _8574_/A sky130_fd_sc_hd__clkbuf_2
X_6537_ _6541_/B _6537_/B vssd1 vssd1 vccd1 vccd1 _6538_/B sky130_fd_sc_hd__and2_1
X_4798_ _4758_/A _4749_/A _4878_/A vssd1 vssd1 vccd1 vccd1 _4799_/D sky130_fd_sc_hd__o21a_1
X_6468_ _8641_/Q _8640_/Q _6468_/C _8644_/Q vssd1 vssd1 vccd1 vccd1 _6471_/B sky130_fd_sc_hd__and4_1
X_6399_ input2/X _8566_/S vssd1 vssd1 vccd1 vccd1 _6464_/B sky130_fd_sc_hd__and2_2
X_8207_ _8325_/A _8229_/B _8323_/C vssd1 vssd1 vccd1 vccd1 _8442_/A sky130_fd_sc_hd__o21ba_1
X_5419_ _8661_/Q _5425_/B vssd1 vssd1 vccd1 vccd1 _5423_/B sky130_fd_sc_hd__or2b_1
XFILLER_87_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8138_ _8138_/A _8201_/B vssd1 vssd1 vccd1 vccd1 _8143_/A sky130_fd_sc_hd__xnor2_2
X_8069_ _8069_/A _8069_/B vssd1 vssd1 vccd1 vccd1 _8072_/C sky130_fd_sc_hd__xnor2_1
XFILLER_101_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5770_ _5757_/A _5770_/B vssd1 vssd1 vccd1 vccd1 _5770_/X sky130_fd_sc_hd__and2b_1
X_4721_ _6600_/B vssd1 vssd1 vccd1 vccd1 _6746_/B sky130_fd_sc_hd__clkbuf_2
X_7440_ _7438_/Y _7339_/B _7439_/Y vssd1 vssd1 vccd1 vccd1 _7441_/B sky130_fd_sc_hd__a21oi_1
X_4652_ _5389_/A _4648_/B _4648_/Y _4651_/X vssd1 vssd1 vccd1 vccd1 _8601_/D sky130_fd_sc_hd__o211a_1
X_7371_ _7371_/A _7413_/B vssd1 vssd1 vccd1 vccd1 _7372_/B sky130_fd_sc_hd__xnor2_1
X_4583_ input2/X vssd1 vssd1 vccd1 vccd1 _6503_/A sky130_fd_sc_hd__clkinv_2
X_6322_ _6322_/A _6322_/B vssd1 vssd1 vccd1 vccd1 _6332_/C sky130_fd_sc_hd__nor2_1
Xclkbuf_4_5_0_wb_clk_i clkbuf_4_5_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _8735_/CLK
+ sky130_fd_sc_hd__clkbuf_2
X_6253_ _6253_/A _6253_/B vssd1 vssd1 vccd1 vccd1 _6253_/X sky130_fd_sc_hd__or2_1
X_5204_ _5139_/D _5203_/X _5220_/A vssd1 vssd1 vccd1 vccd1 _5205_/C sky130_fd_sc_hd__o21a_1
XFILLER_69_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6184_ _5910_/B _5962_/B _5961_/A vssd1 vssd1 vccd1 vccd1 _6185_/A sky130_fd_sc_hd__a21oi_1
X_5135_ _5205_/A _5028_/B _5045_/B _5134_/X _4707_/A vssd1 vssd1 vccd1 vccd1 _5135_/X
+ sky130_fd_sc_hd__o32a_1
X_5066_ _5066_/A _5087_/B vssd1 vssd1 vccd1 vccd1 _5193_/B sky130_fd_sc_hd__and2_1
XFILLER_57_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5968_ _5746_/A _5973_/A _5967_/X vssd1 vssd1 vccd1 vccd1 _5969_/B sky130_fd_sc_hd__o21a_1
XFILLER_25_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4919_ _4919_/A vssd1 vssd1 vccd1 vccd1 _4937_/A sky130_fd_sc_hd__clkbuf_2
X_7707_ _7859_/B _7859_/C vssd1 vssd1 vccd1 vccd1 _7955_/A sky130_fd_sc_hd__nand2_1
XFILLER_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8687_ _8689_/CLK _8687_/D vssd1 vssd1 vccd1 vccd1 _8687_/Q sky130_fd_sc_hd__dfxtp_1
X_5899_ _5899_/A _6221_/B vssd1 vssd1 vccd1 vccd1 _5901_/C sky130_fd_sc_hd__xnor2_1
XFILLER_32_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7638_ _7636_/X _7642_/A vssd1 vssd1 vccd1 vccd1 _7639_/B sky130_fd_sc_hd__and2b_1
XFILLER_4_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7569_ _8723_/Q vssd1 vssd1 vccd1 vccd1 _7618_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_4_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8762__29 vssd1 vssd1 vccd1 vccd1 _8762__29/HI _8857_/A sky130_fd_sc_hd__conb_1
XFILLER_73_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6940_ _6940_/A _7046_/A vssd1 vssd1 vccd1 vccd1 _7047_/A sky130_fd_sc_hd__xor2_1
XFILLER_47_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6871_ _7350_/A vssd1 vssd1 vccd1 vccd1 _7213_/B sky130_fd_sc_hd__buf_2
X_8610_ _8703_/CLK _8610_/D vssd1 vssd1 vccd1 vccd1 _8610_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_62_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5822_ _5861_/A _6255_/A vssd1 vssd1 vccd1 vccd1 _5824_/B sky130_fd_sc_hd__xnor2_1
XFILLER_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8541_ _8541_/A _8541_/B vssd1 vssd1 vccd1 vccd1 _8542_/B sky130_fd_sc_hd__nand2_1
X_5753_ _5754_/A _5754_/B _5754_/C vssd1 vssd1 vccd1 vccd1 _5845_/A sky130_fd_sc_hd__a21oi_1
X_4704_ _7695_/B vssd1 vssd1 vccd1 vccd1 _4707_/A sky130_fd_sc_hd__inv_2
X_8472_ _8372_/A _8372_/B _8471_/X vssd1 vssd1 vccd1 vccd1 _8477_/A sky130_fd_sc_hd__a21oi_1
X_5684_ _5685_/A _5685_/B vssd1 vssd1 vccd1 vccd1 _6049_/B sky130_fd_sc_hd__nor2_1
XFILLER_30_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7423_ _7423_/A _7423_/B vssd1 vssd1 vccd1 vccd1 _7424_/B sky130_fd_sc_hd__xnor2_1
X_4635_ _8597_/Q _4637_/C _4612_/B vssd1 vssd1 vccd1 vccd1 _4635_/Y sky130_fd_sc_hd__o21ai_1
X_7354_ _7454_/B _7364_/C _7353_/Y vssd1 vssd1 vccd1 vccd1 _7355_/C sky130_fd_sc_hd__a21oi_1
X_4566_ _4566_/A vssd1 vssd1 vccd1 vccd1 _8882_/A sky130_fd_sc_hd__clkbuf_1
X_6305_ _6305_/A _6305_/B vssd1 vssd1 vccd1 vccd1 _6320_/B sky130_fd_sc_hd__nor2_1
XFILLER_103_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4497_ _4861_/B vssd1 vssd1 vccd1 vccd1 _4864_/A sky130_fd_sc_hd__clkbuf_1
X_7285_ _7272_/A _7272_/B _7283_/B _7284_/X vssd1 vssd1 vccd1 vccd1 _7473_/B sky130_fd_sc_hd__a31o_1
X_6236_ _6236_/A _6236_/B vssd1 vssd1 vccd1 vccd1 _6236_/Y sky130_fd_sc_hd__nand2_1
XFILLER_69_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6167_ _5978_/A _5978_/B _5979_/B _5979_/A vssd1 vssd1 vccd1 vccd1 _6286_/B sky130_fd_sc_hd__a2bb2o_2
X_5118_ _5237_/B _5118_/B vssd1 vssd1 vccd1 vccd1 _5118_/Y sky130_fd_sc_hd__nand2_1
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6098_ _6095_/Y _6122_/A _6098_/S vssd1 vssd1 vccd1 vccd1 _6099_/C sky130_fd_sc_hd__mux2_1
X_5049_ _5230_/A _5086_/B vssd1 vssd1 vccd1 vccd1 _5200_/C sky130_fd_sc_hd__or2_2
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8807__74 vssd1 vssd1 vccd1 vccd1 _8807__74/HI _8916_/A sky130_fd_sc_hd__conb_1
XFILLER_76_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4420_ _4432_/A vssd1 vssd1 vccd1 vccd1 _4425_/A sky130_fd_sc_hd__buf_2
X_4351_ _4351_/A vssd1 vssd1 vccd1 vccd1 _4351_/Y sky130_fd_sc_hd__inv_2
X_7070_ _7145_/A _6837_/X _7072_/A vssd1 vssd1 vccd1 vccd1 _7147_/A sky130_fd_sc_hd__o21ba_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6021_ _6118_/A _6108_/A _6020_/Y vssd1 vssd1 vccd1 vccd1 _6069_/B sky130_fd_sc_hd__a21oi_1
XFILLER_67_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7972_ _7972_/A _8123_/S vssd1 vssd1 vccd1 vccd1 _7973_/B sky130_fd_sc_hd__xor2_1
X_6923_ _7409_/B _6859_/A _6857_/Y _6862_/A vssd1 vssd1 vccd1 vccd1 _6941_/A sky130_fd_sc_hd__o31ai_2
XFILLER_81_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6854_ _6932_/A _6854_/B vssd1 vssd1 vccd1 vccd1 _6926_/B sky130_fd_sc_hd__xnor2_2
X_6785_ _6785_/A _6785_/B vssd1 vssd1 vccd1 vccd1 _6786_/B sky130_fd_sc_hd__xnor2_1
XFILLER_13_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5805_ _5806_/A _5806_/B _6209_/A vssd1 vssd1 vccd1 vccd1 _5868_/A sky130_fd_sc_hd__a21o_1
XFILLER_22_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5736_ _6174_/A vssd1 vssd1 vccd1 vccd1 _5816_/A sky130_fd_sc_hd__inv_2
X_8524_ _8523_/B _8524_/B vssd1 vssd1 vccd1 vccd1 _8525_/D sky130_fd_sc_hd__and2b_1
X_5667_ _6193_/A _5729_/B _5663_/A _5663_/B _5666_/Y vssd1 vssd1 vccd1 vccd1 _5669_/B
+ sky130_fd_sc_hd__o41a_1
X_8455_ _8066_/A _8166_/X _8370_/B _8367_/Y _8072_/A vssd1 vssd1 vccd1 vccd1 _8464_/A
+ sky130_fd_sc_hd__a32o_1
X_7406_ _7321_/B _7406_/B vssd1 vssd1 vccd1 vccd1 _7406_/X sky130_fd_sc_hd__and2b_1
X_4618_ _8591_/Q _4619_/C _4617_/Y vssd1 vssd1 vccd1 vccd1 _8591_/D sky130_fd_sc_hd__a21oi_1
X_8386_ _8460_/A _8386_/B vssd1 vssd1 vccd1 vccd1 _8394_/A sky130_fd_sc_hd__nor2_1
X_5598_ _5587_/A _5638_/B _5594_/B _5589_/X vssd1 vssd1 vccd1 vccd1 _5661_/B sky130_fd_sc_hd__a211o_1
X_7337_ _7337_/A _7337_/B vssd1 vssd1 vccd1 vccd1 _7338_/B sky130_fd_sc_hd__xor2_2
X_4549_ _4549_/A vssd1 vssd1 vccd1 vccd1 _8878_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_104_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7268_ _7335_/A _7069_/A _7239_/X vssd1 vssd1 vccd1 vccd1 _7269_/A sky130_fd_sc_hd__a21o_1
XFILLER_104_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6219_ _5569_/X _6218_/Y _6219_/S vssd1 vssd1 vccd1 vccd1 _6220_/B sky130_fd_sc_hd__mux2_1
X_7199_ _7198_/A _7198_/B _7203_/A _7203_/B vssd1 vssd1 vccd1 vccd1 _7201_/B sky130_fd_sc_hd__o2bb2a_1
XINSDIODE2_10 _6598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6570_ _8699_/Q _6570_/B vssd1 vssd1 vccd1 vccd1 _6570_/X sky130_fd_sc_hd__and2b_1
X_5521_ _5874_/A _5521_/B _5521_/C _5559_/A vssd1 vssd1 vccd1 vccd1 _5559_/B sky130_fd_sc_hd__nand4_1
X_8240_ _8240_/A _8240_/B vssd1 vssd1 vccd1 vccd1 _8274_/B sky130_fd_sc_hd__xnor2_1
X_5452_ _5540_/A _6316_/A _5451_/X vssd1 vssd1 vccd1 vccd1 _5480_/B sky130_fd_sc_hd__a21o_4
X_4403_ _4406_/A vssd1 vssd1 vccd1 vccd1 _4403_/Y sky130_fd_sc_hd__inv_2
X_8171_ _8473_/S _8196_/A vssd1 vssd1 vccd1 vccd1 _8172_/C sky130_fd_sc_hd__nor2_1
X_5383_ _8658_/Q vssd1 vssd1 vccd1 vccd1 _5400_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7122_ _7120_/A _7120_/B _7121_/X vssd1 vssd1 vccd1 vccd1 _7395_/B sky130_fd_sc_hd__a21oi_1
X_4334_ _4338_/A vssd1 vssd1 vccd1 vccd1 _4334_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7053_ _7392_/A _7053_/B vssd1 vssd1 vccd1 vccd1 _7395_/A sky130_fd_sc_hd__xnor2_2
XFILLER_5_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6004_ _6004_/A _6215_/B vssd1 vssd1 vccd1 vccd1 _6005_/B sky130_fd_sc_hd__xnor2_1
XFILLER_101_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8798__65 vssd1 vssd1 vccd1 vccd1 _8798__65/HI _8907_/A sky130_fd_sc_hd__conb_1
XFILLER_67_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7955_ _7955_/A _8330_/A _7955_/C _7955_/D vssd1 vssd1 vccd1 vccd1 _8026_/A sky130_fd_sc_hd__or4_2
X_6906_ _6711_/A _7102_/B _6785_/B _6905_/X vssd1 vssd1 vccd1 vccd1 _6919_/A sky130_fd_sc_hd__o31a_1
X_7886_ _7886_/A _7960_/B _7886_/C vssd1 vssd1 vccd1 vccd1 _7891_/B sky130_fd_sc_hd__and3_1
X_6837_ _7063_/B _7165_/B vssd1 vssd1 vccd1 vccd1 _6837_/X sky130_fd_sc_hd__and2b_1
XFILLER_50_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6768_ _6768_/A _6768_/B vssd1 vssd1 vccd1 vccd1 _6789_/A sky130_fd_sc_hd__nand2_1
X_8507_ _8506_/B _8506_/C _8506_/A vssd1 vssd1 vccd1 vccd1 _8508_/B sky130_fd_sc_hd__a21oi_1
X_6699_ _6699_/A vssd1 vssd1 vccd1 vccd1 _7169_/A sky130_fd_sc_hd__clkbuf_1
X_5719_ _5806_/B _5719_/B vssd1 vssd1 vccd1 vccd1 _5720_/B sky130_fd_sc_hd__nand2_1
X_8438_ _8425_/A _8425_/B _8437_/Y vssd1 vssd1 vccd1 vccd1 _8486_/A sky130_fd_sc_hd__o21ai_1
X_8369_ _8367_/Y _8306_/B _8368_/Y vssd1 vssd1 vccd1 vccd1 _8371_/A sky130_fd_sc_hd__a21oi_1
X_8738__5 vssd1 vssd1 vccd1 vccd1 _8738__5/HI _8833_/A sky130_fd_sc_hd__conb_1
XFILLER_2_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4952_ _5192_/A _4965_/B _4946_/X _4970_/B _4951_/X vssd1 vssd1 vccd1 vccd1 _4953_/D
+ sky130_fd_sc_hd__o32a_1
X_7740_ _7642_/A _7642_/B _7644_/X _7651_/X _7645_/A vssd1 vssd1 vccd1 vccd1 _7741_/B
+ sky130_fd_sc_hd__a311o_1
X_4883_ _5111_/A _4882_/X vssd1 vssd1 vccd1 vccd1 _5107_/A sky130_fd_sc_hd__or2b_1
X_7671_ _7736_/A _7671_/B vssd1 vssd1 vccd1 vccd1 _7725_/B sky130_fd_sc_hd__xnor2_1
X_6622_ _7465_/A _7434_/B _6619_/Y vssd1 vssd1 vccd1 vccd1 _7293_/A sky130_fd_sc_hd__o21ai_4
XFILLER_20_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6553_ _8710_/Q _6553_/B vssd1 vssd1 vccd1 vccd1 _6553_/X sky130_fd_sc_hd__and2b_1
XFILLER_9_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6484_ _6479_/X _6481_/X _7540_/A _7546_/A vssd1 vssd1 vccd1 vccd1 _6484_/X sky130_fd_sc_hd__a211o_1
X_5504_ _5792_/B _5780_/B _5780_/C vssd1 vssd1 vccd1 vccd1 _5896_/A sky130_fd_sc_hd__nand3_4
X_5435_ _4581_/B _5434_/C _5634_/A vssd1 vssd1 vccd1 vccd1 _5436_/C sky130_fd_sc_hd__o21ai_1
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8223_ _8223_/A _8223_/B vssd1 vssd1 vccd1 vccd1 _8235_/A sky130_fd_sc_hd__xnor2_1
XFILLER_87_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8154_ _8155_/A _8390_/A vssd1 vssd1 vccd1 vccd1 _8200_/A sky130_fd_sc_hd__nand2_1
X_5366_ _8674_/Q vssd1 vssd1 vccd1 vccd1 _5374_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_99_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5297_ _5323_/A vssd1 vssd1 vccd1 vccd1 _5359_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7105_ _7105_/A _7105_/B _7105_/C vssd1 vssd1 vccd1 vccd1 _7125_/C sky130_fd_sc_hd__and3_1
X_8085_ _8243_/B _8085_/B vssd1 vssd1 vccd1 vccd1 _8087_/A sky130_fd_sc_hd__or2_1
X_7036_ _7036_/A _7036_/B vssd1 vssd1 vccd1 vccd1 _7304_/A sky130_fd_sc_hd__xnor2_1
XFILLER_87_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7938_ _7938_/A _7938_/B vssd1 vssd1 vccd1 vccd1 _7940_/C sky130_fd_sc_hd__or2_1
XFILLER_35_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7869_ _7869_/A _7869_/B vssd1 vssd1 vccd1 vccd1 _8330_/A sky130_fd_sc_hd__xnor2_4
XFILLER_23_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5220_ _5220_/A _5220_/B _5220_/C _5220_/D vssd1 vssd1 vccd1 vccd1 _5220_/X sky130_fd_sc_hd__or4_1
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5151_ _4661_/A _5028_/C _4916_/A vssd1 vssd1 vccd1 vccd1 _5151_/X sky130_fd_sc_hd__o21a_1
XFILLER_96_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5082_ _5044_/B _5143_/B _5065_/X _5081_/X _4711_/B vssd1 vssd1 vccd1 vccd1 _5082_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_69_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8910_ _8910_/A _4421_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[9] sky130_fd_sc_hd__ebufn_8
X_8768__35 vssd1 vssd1 vccd1 vccd1 _8768__35/HI _8863_/A sky130_fd_sc_hd__conb_1
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8841_ _8841_/A _4344_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[10] sky130_fd_sc_hd__ebufn_8
XFILLER_64_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7723_ _7836_/A vssd1 vssd1 vccd1 vccd1 _8054_/A sky130_fd_sc_hd__clkbuf_2
X_5984_ _5891_/A _5982_/X _5983_/X vssd1 vssd1 vccd1 vccd1 _6191_/A sky130_fd_sc_hd__a21o_1
X_4935_ _5244_/B vssd1 vssd1 vccd1 vccd1 _5207_/B sky130_fd_sc_hd__clkbuf_2
X_4866_ _4795_/C _4899_/C _4822_/A vssd1 vssd1 vccd1 vccd1 _4867_/B sky130_fd_sc_hd__a21oi_1
XFILLER_32_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7654_ _7654_/A _7654_/B vssd1 vssd1 vccd1 vccd1 _8145_/A sky130_fd_sc_hd__xnor2_4
X_6605_ _7540_/A _6605_/B vssd1 vssd1 vccd1 vccd1 _6605_/X sky130_fd_sc_hd__and2b_1
X_4797_ _4828_/A _4839_/B _4834_/C _4847_/A vssd1 vssd1 vccd1 vccd1 _4878_/A sky130_fd_sc_hd__or4b_2
X_7585_ _8566_/S vssd1 vssd1 vccd1 vccd1 _8543_/S sky130_fd_sc_hd__buf_2
X_6536_ _6536_/A _6536_/B vssd1 vssd1 vccd1 vccd1 _6537_/B sky130_fd_sc_hd__or2_1
XFILLER_21_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6467_ _8647_/Q _8646_/Q _8654_/Q _6467_/D vssd1 vssd1 vccd1 vccd1 _6472_/C sky130_fd_sc_hd__nor4_1
X_6398_ _6403_/B _7555_/A vssd1 vssd1 vccd1 vccd1 _8566_/S sky130_fd_sc_hd__or2_4
X_8206_ _8206_/A _8229_/B vssd1 vssd1 vccd1 vccd1 _8323_/C sky130_fd_sc_hd__and2_1
X_5418_ _5425_/B _5432_/A vssd1 vssd1 vccd1 vccd1 _5427_/A sky130_fd_sc_hd__or2b_1
XFILLER_99_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5349_ _8649_/Q _5351_/C _5323_/X vssd1 vssd1 vccd1 vccd1 _5350_/B sky130_fd_sc_hd__o21ai_1
X_8137_ _8137_/A _8137_/B vssd1 vssd1 vccd1 vccd1 _8201_/B sky130_fd_sc_hd__xnor2_1
XFILLER_101_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8068_ _8167_/A _8291_/A _8067_/Y vssd1 vssd1 vccd1 vccd1 _8069_/B sky130_fd_sc_hd__o21a_1
X_7019_ _7018_/A _7018_/B _7018_/C vssd1 vssd1 vccd1 vccd1 _7019_/X sky130_fd_sc_hd__o21a_1
XFILLER_46_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4720_ _4720_/A vssd1 vssd1 vccd1 vccd1 _6600_/B sky130_fd_sc_hd__inv_2
X_4651_ _8567_/A vssd1 vssd1 vccd1 vccd1 _4651_/X sky130_fd_sc_hd__buf_2
X_7370_ _7370_/A _7454_/C vssd1 vssd1 vccd1 vccd1 _7413_/B sky130_fd_sc_hd__xor2_1
X_4582_ _8581_/Q _4582_/B vssd1 vssd1 vccd1 vccd1 _8581_/D sky130_fd_sc_hd__nor2_1
XFILLER_6_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6321_ _6321_/A _6321_/B vssd1 vssd1 vccd1 vccd1 _6322_/B sky130_fd_sc_hd__and2_1
X_6252_ _6224_/A _6224_/B _6227_/A vssd1 vssd1 vccd1 vccd1 _6260_/A sky130_fd_sc_hd__a21oi_1
X_5203_ _4923_/A _5231_/B _5109_/C _5202_/X vssd1 vssd1 vccd1 vccd1 _5203_/X sky130_fd_sc_hd__o31a_1
X_6183_ _6286_/B _6183_/B vssd1 vssd1 vccd1 vccd1 _6186_/A sky130_fd_sc_hd__xnor2_4
X_5134_ _5164_/C _5127_/X _5128_/X _5166_/A _5133_/X vssd1 vssd1 vccd1 vccd1 _5134_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_69_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5065_ _5065_/A _5155_/B _5179_/B _5065_/D vssd1 vssd1 vccd1 vccd1 _5065_/X sky130_fd_sc_hd__or4_1
XFILLER_16_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5967_ _5967_/A _6273_/S vssd1 vssd1 vccd1 vccd1 _5967_/X sky130_fd_sc_hd__or2_1
X_8686_ _8689_/CLK _8686_/D vssd1 vssd1 vccd1 vccd1 _8686_/Q sky130_fd_sc_hd__dfxtp_1
X_4918_ _5127_/A vssd1 vssd1 vccd1 vccd1 _5166_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_52_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7706_ _7713_/A _7713_/B vssd1 vssd1 vccd1 vccd1 _7859_/C sky130_fd_sc_hd__xor2_2
X_5898_ _6002_/A vssd1 vssd1 vccd1 vccd1 _6221_/B sky130_fd_sc_hd__inv_2
XFILLER_32_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7637_ _8617_/Q _7596_/B vssd1 vssd1 vccd1 vccd1 _7642_/A sky130_fd_sc_hd__or2b_2
X_4849_ _4937_/B _4849_/B vssd1 vssd1 vccd1 vccd1 _4977_/A sky130_fd_sc_hd__nor2_1
XFILLER_20_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7568_ _7618_/B vssd1 vssd1 vccd1 vccd1 _7617_/B sky130_fd_sc_hd__clkbuf_2
X_6519_ _6515_/A _5362_/X _6508_/X _6518_/X vssd1 vssd1 vccd1 vccd1 _8700_/D sky130_fd_sc_hd__a22o_1
X_7499_ _7499_/A vssd1 vssd1 vccd1 vccd1 _7499_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6870_ _6870_/A _6870_/B vssd1 vssd1 vccd1 vccd1 _7350_/A sky130_fd_sc_hd__nand2_2
XFILLER_19_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5821_ _5821_/A vssd1 vssd1 vccd1 vccd1 _6255_/A sky130_fd_sc_hd__buf_2
XFILLER_22_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5752_ _5810_/A _5752_/B vssd1 vssd1 vccd1 vccd1 _5754_/C sky130_fd_sc_hd__or2_1
X_8540_ _8540_/A _8716_/Q vssd1 vssd1 vccd1 vccd1 _8541_/B sky130_fd_sc_hd__or2b_1
X_4703_ _6553_/B _7695_/B _5226_/A vssd1 vssd1 vccd1 vccd1 _5029_/A sky130_fd_sc_hd__and3_1
X_8471_ _8371_/A _8471_/B vssd1 vssd1 vccd1 vccd1 _8471_/X sky130_fd_sc_hd__and2b_1
X_5683_ _5952_/A _5943_/A _6037_/B _5673_/A _6193_/A vssd1 vssd1 vccd1 vccd1 _5685_/B
+ sky130_fd_sc_hd__o32a_1
X_7422_ _7422_/A _7422_/B vssd1 vssd1 vccd1 vccd1 _7423_/B sky130_fd_sc_hd__xnor2_1
X_4634_ _4637_/C _4634_/B vssd1 vssd1 vccd1 vccd1 _8596_/D sky130_fd_sc_hd__nor2_1
X_7353_ _6892_/B _6958_/B _7352_/X vssd1 vssd1 vccd1 vccd1 _7353_/Y sky130_fd_sc_hd__o21ai_1
X_4565_ _8628_/Q _4567_/B vssd1 vssd1 vccd1 vccd1 _4566_/A sky130_fd_sc_hd__and2_1
X_6304_ _6306_/A _6306_/B _6094_/A vssd1 vssd1 vccd1 vccd1 _6305_/B sky130_fd_sc_hd__a21o_1
X_7284_ _7469_/B _7469_/A vssd1 vssd1 vccd1 vccd1 _7284_/X sky130_fd_sc_hd__and2b_1
X_4496_ _7643_/B vssd1 vssd1 vccd1 vccd1 _4861_/B sky130_fd_sc_hd__buf_2
XFILLER_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6235_ _6236_/A _6235_/B vssd1 vssd1 vccd1 vccd1 _6312_/B sky130_fd_sc_hd__xnor2_1
XFILLER_103_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6166_ _6011_/A _6011_/B _6165_/X vssd1 vssd1 vccd1 vccd1 _6232_/A sky130_fd_sc_hd__a21o_1
XFILLER_84_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5117_ _5127_/A _5220_/B _5212_/B vssd1 vssd1 vccd1 vccd1 _5118_/B sky130_fd_sc_hd__nor3_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6097_ _6120_/A _6097_/B vssd1 vssd1 vccd1 vccd1 _6098_/S sky130_fd_sc_hd__nand2_1
X_5048_ _5199_/C _5209_/C vssd1 vssd1 vccd1 vccd1 _5086_/B sky130_fd_sc_hd__or2_1
XFILLER_72_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6999_ _6999_/A _7000_/B vssd1 vssd1 vccd1 vccd1 _7328_/A sky130_fd_sc_hd__nor2_1
XFILLER_21_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8669_ _8674_/CLK _8669_/D vssd1 vssd1 vccd1 vccd1 _8669_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_21_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8822__89 vssd1 vssd1 vccd1 vccd1 _8822__89/HI _8931_/A sky130_fd_sc_hd__conb_1
XFILLER_75_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4350_ _4351_/A vssd1 vssd1 vccd1 vccd1 _4350_/Y sky130_fd_sc_hd__inv_2
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6020_ _6020_/A _6020_/B vssd1 vssd1 vccd1 vccd1 _6020_/Y sky130_fd_sc_hd__nand2_2
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7971_ _7878_/A _8410_/A _7880_/B _7880_/A vssd1 vssd1 vccd1 vccd1 _8045_/A sky130_fd_sc_hd__a22o_1
X_6922_ _6948_/A _6948_/B vssd1 vssd1 vccd1 vccd1 _6949_/A sky130_fd_sc_hd__xnor2_1
XFILLER_54_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6853_ _6853_/A _7432_/A vssd1 vssd1 vccd1 vccd1 _6854_/B sky130_fd_sc_hd__xnor2_2
XFILLER_62_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5804_ _5713_/X _5788_/B _5981_/B vssd1 vssd1 vccd1 vccd1 _6209_/A sky130_fd_sc_hd__o21ai_4
X_6784_ _6784_/A _6784_/B vssd1 vssd1 vccd1 vccd1 _6785_/B sky130_fd_sc_hd__xnor2_1
XFILLER_50_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5735_ _5859_/B _5944_/B vssd1 vssd1 vccd1 vccd1 _6174_/A sky130_fd_sc_hd__nand2_2
XFILLER_13_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8523_ _8524_/B _8523_/B vssd1 vssd1 vccd1 vccd1 _8529_/B sky130_fd_sc_hd__and2b_1
X_5666_ _6193_/A _5747_/B _5729_/B vssd1 vssd1 vccd1 vccd1 _5666_/Y sky130_fd_sc_hd__o21ai_1
X_8454_ _8454_/A _8454_/B vssd1 vssd1 vccd1 vccd1 _8465_/A sky130_fd_sc_hd__xnor2_1
X_7405_ _7405_/A _7405_/B vssd1 vssd1 vccd1 vccd1 _7425_/A sky130_fd_sc_hd__xnor2_1
X_4617_ _8591_/Q _4619_/C _4607_/X vssd1 vssd1 vccd1 vccd1 _4617_/Y sky130_fd_sc_hd__o21ai_1
X_8385_ _8383_/Y _8349_/B _8384_/Y vssd1 vssd1 vccd1 vccd1 _8422_/A sky130_fd_sc_hd__a21o_1
X_5597_ _7643_/B _8660_/Q vssd1 vssd1 vccd1 vccd1 _5660_/A sky130_fd_sc_hd__or2b_1
XFILLER_104_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7336_ _7280_/A _7102_/A _7336_/S vssd1 vssd1 vccd1 vccd1 _7337_/B sky130_fd_sc_hd__mux2_1
XFILLER_89_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4548_ _8624_/Q _4552_/B vssd1 vssd1 vccd1 vccd1 _4549_/A sky130_fd_sc_hd__and2_1
X_4479_ _6605_/B _6603_/B _4479_/C _4478_/X vssd1 vssd1 vccd1 vccd1 _4541_/A sky130_fd_sc_hd__or4b_1
X_7267_ _7267_/A _7267_/B vssd1 vssd1 vccd1 vccd1 _7272_/A sky130_fd_sc_hd__xor2_1
XFILLER_77_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6218_ _6218_/A _6218_/B vssd1 vssd1 vccd1 vccd1 _6218_/Y sky130_fd_sc_hd__nor2_1
X_7198_ _7198_/A _7198_/B vssd1 vssd1 vccd1 vccd1 _7203_/B sky130_fd_sc_hd__xnor2_1
XFILLER_58_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_11 _7060_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6149_ _6151_/A _6154_/D vssd1 vssd1 vccd1 vccd1 _6150_/B sky130_fd_sc_hd__xor2_1
XFILLER_38_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5520_ _5566_/A _5784_/A _5525_/A vssd1 vssd1 vccd1 vccd1 _5559_/A sky130_fd_sc_hd__or3_1
XFILLER_8_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5451_ _8669_/Q _8606_/Q vssd1 vssd1 vccd1 vccd1 _5451_/X sky130_fd_sc_hd__and2b_1
X_4402_ _4406_/A vssd1 vssd1 vccd1 vccd1 _4402_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8170_ _8368_/A vssd1 vssd1 vccd1 vccd1 _8473_/S sky130_fd_sc_hd__dlymetal6s2s_1
X_5382_ _8659_/Q vssd1 vssd1 vccd1 vccd1 _5404_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_7121_ _7392_/A _7293_/B vssd1 vssd1 vccd1 vccd1 _7121_/X sky130_fd_sc_hd__and2_1
X_4333_ _4464_/A vssd1 vssd1 vccd1 vccd1 _4338_/A sky130_fd_sc_hd__clkbuf_2
X_7052_ _7050_/Y _7052_/B vssd1 vssd1 vccd1 vccd1 _7053_/B sky130_fd_sc_hd__and2b_1
XFILLER_59_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6003_ _5899_/A _6002_/A _5901_/A vssd1 vssd1 vccd1 vccd1 _6215_/B sky130_fd_sc_hd__a21oi_1
XFILLER_39_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7954_ _8208_/A _8118_/B _8118_/C _7859_/C _7950_/A vssd1 vssd1 vccd1 vccd1 _7956_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_27_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6905_ _6905_/A _6786_/B vssd1 vssd1 vccd1 vccd1 _6905_/X sky130_fd_sc_hd__or2b_1
XFILLER_82_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7885_ _7885_/A _7972_/A vssd1 vssd1 vccd1 vccd1 _7891_/A sky130_fd_sc_hd__nor2_1
XFILLER_24_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6836_ _6836_/A _6836_/B vssd1 vssd1 vccd1 vccd1 _7165_/B sky130_fd_sc_hd__xnor2_4
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6767_ _7109_/A _7109_/B _6766_/X vssd1 vssd1 vccd1 vccd1 _6865_/B sky130_fd_sc_hd__o21ai_1
XFILLER_10_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5718_ _5718_/A _5718_/B vssd1 vssd1 vccd1 vccd1 _5719_/B sky130_fd_sc_hd__or2_1
X_8506_ _8506_/A _8506_/B _8506_/C vssd1 vssd1 vccd1 vccd1 _8508_/A sky130_fd_sc_hd__and3_1
X_6698_ _6697_/A _6697_/B _6697_/C vssd1 vssd1 vccd1 vccd1 _6704_/B sky130_fd_sc_hd__a21o_1
X_5649_ _5859_/B vssd1 vssd1 vccd1 vccd1 _6097_/B sky130_fd_sc_hd__clkbuf_2
X_8437_ _8437_/A _8437_/B vssd1 vssd1 vccd1 vccd1 _8437_/Y sky130_fd_sc_hd__nand2_1
X_8368_ _8368_/A _8368_/B vssd1 vssd1 vccd1 vccd1 _8368_/Y sky130_fd_sc_hd__nor2_1
XFILLER_104_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7319_ _7401_/B _7319_/B vssd1 vssd1 vccd1 vccd1 _7320_/B sky130_fd_sc_hd__xnor2_1
XFILLER_49_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8299_ _8299_/A _8299_/B vssd1 vssd1 vccd1 vccd1 _8351_/A sky130_fd_sc_hd__xor2_1
XFILLER_49_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4951_ _5240_/B _5126_/B _4987_/B _5223_/D vssd1 vssd1 vccd1 vccd1 _4951_/X sky130_fd_sc_hd__or4_1
XFILLER_17_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4882_ _4885_/B _4890_/B vssd1 vssd1 vccd1 vccd1 _4882_/X sky130_fd_sc_hd__or2_1
X_7670_ _7661_/C _7663_/Y _7670_/S vssd1 vssd1 vccd1 vccd1 _7671_/B sky130_fd_sc_hd__mux2_1
XFILLER_32_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6621_ _6916_/A vssd1 vssd1 vccd1 vccd1 _7434_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_20_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6552_ _8710_/Q _6553_/B vssd1 vssd1 vccd1 vccd1 _6582_/B sky130_fd_sc_hd__xnor2_2
X_6483_ _8713_/Q vssd1 vssd1 vccd1 vccd1 _7546_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5503_ _5503_/A vssd1 vssd1 vccd1 vccd1 _5792_/B sky130_fd_sc_hd__clkbuf_2
X_5434_ _5634_/A _5434_/B _5434_/C vssd1 vssd1 vccd1 vccd1 _5436_/B sky130_fd_sc_hd__or3_1
X_8222_ _8319_/A _8319_/B vssd1 vssd1 vccd1 vccd1 _8223_/B sky130_fd_sc_hd__xnor2_1
X_8153_ _8054_/A _7836_/C _8365_/B vssd1 vssd1 vccd1 vccd1 _8390_/A sky130_fd_sc_hd__o21a_2
XFILLER_99_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7104_ _7124_/D _7124_/C _7127_/B _7107_/A vssd1 vssd1 vccd1 vccd1 _7125_/B sky130_fd_sc_hd__o2bb2a_1
X_5365_ _6353_/B vssd1 vssd1 vccd1 vccd1 _6368_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_5296_ _5296_/A _6502_/A vssd1 vssd1 vccd1 vccd1 _5323_/A sky130_fd_sc_hd__and2_1
XFILLER_59_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8084_ _8084_/A _8002_/B vssd1 vssd1 vccd1 vccd1 _8094_/A sky130_fd_sc_hd__or2b_1
XFILLER_101_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7035_ _7317_/A _7317_/B vssd1 vssd1 vccd1 vccd1 _7036_/B sky130_fd_sc_hd__xnor2_1
XFILLER_19_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7937_ _7936_/A _7936_/B _7936_/C vssd1 vssd1 vccd1 vccd1 _7938_/B sky130_fd_sc_hd__o21a_1
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7868_ _7867_/B _7867_/C _7867_/A vssd1 vssd1 vccd1 vccd1 _7881_/B sky130_fd_sc_hd__a21o_1
X_8740__7 vssd1 vssd1 vccd1 vccd1 _8740__7/HI _8835_/A sky130_fd_sc_hd__conb_1
Xclkbuf_2_0_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
X_6819_ _6819_/A _6819_/B vssd1 vssd1 vccd1 vccd1 _6820_/B sky130_fd_sc_hd__xnor2_1
XFILLER_11_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7799_ _7748_/A _7748_/B _7798_/X vssd1 vssd1 vccd1 vccd1 _7901_/A sky130_fd_sc_hd__a21oi_2
XFILLER_51_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5150_ _5194_/C _5022_/B _5131_/A _4960_/A vssd1 vssd1 vccd1 vccd1 _5150_/X sky130_fd_sc_hd__o31a_1
XFILLER_69_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5081_ _5073_/X _5078_/X _5080_/Y vssd1 vssd1 vccd1 vccd1 _5081_/X sky130_fd_sc_hd__a21o_1
XFILLER_84_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8840_ _8840_/A _4343_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[9] sky130_fd_sc_hd__ebufn_8
XFILLER_37_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5983_ _5983_/A _5983_/B vssd1 vssd1 vccd1 vccd1 _5983_/X sky130_fd_sc_hd__and2_1
X_4934_ _5087_/A _4820_/X _5007_/A vssd1 vssd1 vccd1 vccd1 _4987_/B sky130_fd_sc_hd__a21o_1
X_7722_ _7722_/A _7722_/B vssd1 vssd1 vccd1 vccd1 _7836_/A sky130_fd_sc_hd__nand2_1
X_4865_ _4903_/B _4827_/A _5066_/A _4864_/X vssd1 vssd1 vccd1 vccd1 _5185_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_20_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7653_ _7651_/X _7741_/A vssd1 vssd1 vccd1 vccd1 _7654_/B sky130_fd_sc_hd__and2b_1
X_6604_ _6745_/A _6747_/A _6745_/B _6602_/Y _6811_/B vssd1 vssd1 vccd1 vccd1 _6826_/B
+ sky130_fd_sc_hd__a311o_1
X_4796_ _4823_/B _4796_/B vssd1 vssd1 vccd1 vccd1 _4899_/B sky130_fd_sc_hd__or2_2
X_7584_ _8578_/A vssd1 vssd1 vccd1 vccd1 _7584_/X sky130_fd_sc_hd__clkbuf_2
X_6535_ _6536_/A _6536_/B vssd1 vssd1 vccd1 vccd1 _6541_/B sky130_fd_sc_hd__nand2_1
XFILLER_21_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6466_ _8639_/Q _6466_/B _8643_/Q _6466_/D vssd1 vssd1 vccd1 vccd1 _6467_/D sky130_fd_sc_hd__or4_1
X_8205_ _8205_/A _8450_/A vssd1 vssd1 vccd1 vccd1 _8229_/B sky130_fd_sc_hd__nor2_1
X_6397_ _6397_/A _6397_/B _6397_/C vssd1 vssd1 vccd1 vccd1 _7555_/A sky130_fd_sc_hd__and3_4
X_5417_ _5411_/B _5410_/X _5415_/Y _5416_/X _4746_/X vssd1 vssd1 vccd1 vccd1 _8660_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_99_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5348_ _8649_/Q _5351_/C vssd1 vssd1 vccd1 vccd1 _5350_/A sky130_fd_sc_hd__and2_1
X_8136_ _8211_/B _8136_/B vssd1 vssd1 vccd1 vccd1 _8137_/B sky130_fd_sc_hd__nor2_1
XFILLER_99_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8067_ _8196_/A _8370_/A vssd1 vssd1 vccd1 vccd1 _8067_/Y sky130_fd_sc_hd__nand2_1
X_7018_ _7018_/A _7018_/B _7018_/C vssd1 vssd1 vccd1 vccd1 _7018_/Y sky130_fd_sc_hd__nor3_1
XFILLER_87_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5279_ _8567_/A vssd1 vssd1 vccd1 vccd1 _5279_/X sky130_fd_sc_hd__buf_2
XFILLER_28_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4650_ _5296_/A vssd1 vssd1 vccd1 vccd1 _8567_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6320_ _6320_/A _6320_/B _6320_/C vssd1 vssd1 vccd1 vccd1 _6320_/X sky130_fd_sc_hd__or3_1
X_4581_ _8531_/A _4581_/B vssd1 vssd1 vccd1 vccd1 _4582_/B sky130_fd_sc_hd__nand2_1
X_6251_ _6251_/A _6251_/B vssd1 vssd1 vccd1 vccd1 _6261_/A sky130_fd_sc_hd__xnor2_1
XFILLER_103_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8828__95 vssd1 vssd1 vccd1 vccd1 _8828__95/HI _8937_/A sky130_fd_sc_hd__conb_1
XFILLER_88_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5202_ _5230_/A _5223_/A _5202_/C _5202_/D vssd1 vssd1 vccd1 vccd1 _5202_/X sky130_fd_sc_hd__or4_1
X_6182_ _6182_/A _6182_/B vssd1 vssd1 vccd1 vccd1 _6183_/B sky130_fd_sc_hd__xnor2_2
X_5133_ _5237_/A _5143_/B _5218_/D _5132_/X vssd1 vssd1 vccd1 vccd1 _5133_/X sky130_fd_sc_hd__a211o_1
XFILLER_57_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5064_ _5064_/A _5064_/B _5064_/C vssd1 vssd1 vccd1 vccd1 _5064_/X sky130_fd_sc_hd__or3_1
XFILLER_65_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5966_ _5907_/A _5907_/B _5965_/X vssd1 vssd1 vccd1 vccd1 _6010_/A sky130_fd_sc_hd__a21oi_1
X_8685_ _8695_/CLK _8685_/D vssd1 vssd1 vccd1 vccd1 _8685_/Q sky130_fd_sc_hd__dfxtp_1
X_4917_ _4917_/A vssd1 vssd1 vccd1 vccd1 _4928_/A sky130_fd_sc_hd__inv_2
X_5897_ _6204_/B _6134_/B _5997_/A vssd1 vssd1 vccd1 vccd1 _6002_/A sky130_fd_sc_hd__a21oi_2
XFILLER_40_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7705_ _7712_/A _7712_/B _7681_/A vssd1 vssd1 vccd1 vccd1 _7713_/A sky130_fd_sc_hd__a21o_2
X_4848_ _4848_/A _4848_/B _4848_/C _4839_/A vssd1 vssd1 vccd1 vccd1 _4937_/B sky130_fd_sc_hd__or4b_2
XFILLER_32_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7636_ _8720_/Q _8617_/Q vssd1 vssd1 vccd1 vccd1 _7636_/X sky130_fd_sc_hd__and2b_1
XFILLER_32_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4779_ _4790_/A _4779_/B vssd1 vssd1 vccd1 vccd1 _4779_/Y sky130_fd_sc_hd__nand2_1
X_7567_ _8717_/Q vssd1 vssd1 vccd1 vccd1 _7618_/B sky130_fd_sc_hd__clkbuf_1
X_6518_ _6518_/A _6518_/B vssd1 vssd1 vccd1 vccd1 _6518_/X sky130_fd_sc_hd__xor2_1
X_7498_ _6325_/X _8705_/Q _7492_/X _7497_/X vssd1 vssd1 vccd1 vccd1 _8705_/D sky130_fd_sc_hd__o22a_1
X_6449_ _6449_/A vssd1 vssd1 vccd1 vccd1 _8689_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8119_ _8119_/A _8131_/B vssd1 vssd1 vccd1 vccd1 _8120_/B sky130_fd_sc_hd__xnor2_1
XFILLER_87_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5820_ _5820_/A _5962_/A _6174_/A vssd1 vssd1 vccd1 vccd1 _5821_/A sky130_fd_sc_hd__and3_1
XFILLER_22_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5751_ _5751_/A _5751_/B _5751_/C vssd1 vssd1 vccd1 vccd1 _5752_/B sky130_fd_sc_hd__and3_1
XFILLER_22_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4702_ _4702_/A _4702_/B vssd1 vssd1 vccd1 vccd1 _4716_/A sky130_fd_sc_hd__nor2_1
X_8470_ _8374_/A _8374_/B _8469_/X vssd1 vssd1 vccd1 vccd1 _8478_/A sky130_fd_sc_hd__a21oi_1
X_7421_ _7455_/B _7447_/B _7359_/C _7378_/A vssd1 vssd1 vccd1 vccd1 _7422_/B sky130_fd_sc_hd__a31o_1
X_5682_ _5682_/A _6030_/B vssd1 vssd1 vccd1 vccd1 _6037_/B sky130_fd_sc_hd__xnor2_1
X_4633_ _8596_/Q _4632_/B _4607_/X vssd1 vssd1 vccd1 vccd1 _4634_/B sky130_fd_sc_hd__o21ai_1
XFILLER_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7352_ _7352_/A _7352_/B _7352_/C vssd1 vssd1 vccd1 vccd1 _7352_/X sky130_fd_sc_hd__or3_1
X_4564_ _4564_/A vssd1 vssd1 vccd1 vccd1 _8881_/A sky130_fd_sc_hd__clkbuf_1
X_7283_ _7283_/A _7283_/B vssd1 vssd1 vccd1 vccd1 _7469_/A sky130_fd_sc_hd__xnor2_2
X_6303_ _6303_/A _6303_/B vssd1 vssd1 vccd1 vccd1 _6305_/A sky130_fd_sc_hd__xnor2_1
XFILLER_103_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4495_ _8618_/Q vssd1 vssd1 vccd1 vccd1 _7643_/B sky130_fd_sc_hd__clkbuf_2
X_6234_ _6234_/A _6234_/B vssd1 vssd1 vccd1 vccd1 _6235_/B sky130_fd_sc_hd__xor2_2
XFILLER_97_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6165_ _6010_/A _6165_/B vssd1 vssd1 vccd1 vccd1 _6165_/X sky130_fd_sc_hd__and2b_1
XFILLER_85_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5116_ _5116_/A vssd1 vssd1 vccd1 vccd1 _5212_/B sky130_fd_sc_hd__clkbuf_2
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6096_ _6096_/A _6096_/B vssd1 vssd1 vccd1 vccd1 _6122_/A sky130_fd_sc_hd__nor2_1
X_5047_ _5047_/A _5047_/B vssd1 vssd1 vccd1 vccd1 _5209_/C sky130_fd_sc_hd__nor2_1
XFILLER_27_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6998_ _6883_/A _6883_/B _6882_/B _6997_/Y vssd1 vssd1 vccd1 vccd1 _7306_/A sky130_fd_sc_hd__o2bb2a_1
X_5949_ _5952_/C vssd1 vssd1 vccd1 vccd1 _6119_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_43_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8668_ _8674_/CLK _8668_/D vssd1 vssd1 vccd1 vccd1 _8668_/Q sky130_fd_sc_hd__dfxtp_1
X_8599_ _8600_/CLK _8599_/D vssd1 vssd1 vccd1 vccd1 _8599_/Q sky130_fd_sc_hd__dfxtp_1
X_7619_ _7619_/A _7623_/B vssd1 vssd1 vccd1 vccd1 _7620_/B sky130_fd_sc_hd__nand2_1
XFILLER_4_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7970_ _7970_/A _8044_/A vssd1 vssd1 vccd1 vccd1 _8046_/A sky130_fd_sc_hd__or2_1
X_6921_ _6950_/A _6921_/B vssd1 vssd1 vccd1 vccd1 _6948_/B sky130_fd_sc_hd__xnor2_1
XFILLER_81_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6852_ _7310_/A vssd1 vssd1 vccd1 vccd1 _6932_/A sky130_fd_sc_hd__clkbuf_2
X_5803_ _6020_/A _6218_/A vssd1 vssd1 vccd1 vccd1 _5981_/B sky130_fd_sc_hd__nand2_4
X_6783_ _7348_/B _7352_/B vssd1 vssd1 vccd1 vccd1 _6784_/B sky130_fd_sc_hd__nor2_1
X_8522_ _7499_/X _8517_/X _8520_/X _8521_/Y vssd1 vssd1 vccd1 vccd1 _8725_/D sky130_fd_sc_hd__a31oi_1
XFILLER_13_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5734_ _5941_/B _6273_/S _5841_/A vssd1 vssd1 vccd1 vccd1 _5738_/A sky130_fd_sc_hd__o21a_1
X_5665_ _6030_/B vssd1 vssd1 vccd1 vccd1 _5747_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_8453_ _8453_/A _8453_/B vssd1 vssd1 vccd1 vccd1 _8454_/B sky130_fd_sc_hd__xnor2_1
X_7404_ _6932_/A _6926_/A _7312_/A _7310_/X vssd1 vssd1 vccd1 vccd1 _7405_/B sky130_fd_sc_hd__o22a_1
X_4616_ _4619_/C _4616_/B vssd1 vssd1 vccd1 vccd1 _8590_/D sky130_fd_sc_hd__nor2_1
X_8384_ _8384_/A _8384_/B vssd1 vssd1 vccd1 vccd1 _8384_/Y sky130_fd_sc_hd__nor2_1
X_7335_ _7335_/A _7335_/B vssd1 vssd1 vccd1 vccd1 _7337_/A sky130_fd_sc_hd__nand2_1
X_5596_ _5948_/A vssd1 vssd1 vccd1 vccd1 _5940_/B sky130_fd_sc_hd__inv_2
X_4547_ _4547_/A vssd1 vssd1 vccd1 vccd1 _8877_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4478_ _6596_/B vssd1 vssd1 vccd1 vccd1 _4478_/X sky130_fd_sc_hd__clkbuf_1
X_7266_ _7286_/A _7286_/B _7286_/C vssd1 vssd1 vccd1 vccd1 _7266_/X sky130_fd_sc_hd__a21o_1
X_7197_ _7465_/A _7055_/X _7196_/X vssd1 vssd1 vccd1 vccd1 _7203_/A sky130_fd_sc_hd__o21a_1
X_6217_ _5993_/A _6219_/S _5994_/B _6218_/B vssd1 vssd1 vccd1 vccd1 _6220_/A sky130_fd_sc_hd__a22o_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6148_ _6148_/A _6148_/B vssd1 vssd1 vccd1 vccd1 _6154_/D sky130_fd_sc_hd__xor2_1
XFILLER_97_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_12 _8554_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6079_ _6046_/A _6045_/B _6044_/X vssd1 vssd1 vccd1 vccd1 _6079_/X sky130_fd_sc_hd__o21ba_1
XFILLER_72_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5450_ _5450_/A _5450_/B vssd1 vssd1 vccd1 vccd1 _5480_/A sky130_fd_sc_hd__nor2_4
X_4401_ _4401_/A vssd1 vssd1 vccd1 vccd1 _4406_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5381_ _8661_/Q vssd1 vssd1 vccd1 vccd1 _5432_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4332_ _4456_/A vssd1 vssd1 vccd1 vccd1 _4464_/A sky130_fd_sc_hd__buf_6
X_7120_ _7120_/A _7120_/B vssd1 vssd1 vccd1 vccd1 _7293_/B sky130_fd_sc_hd__xor2_1
XFILLER_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_2_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_5_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
X_7051_ _7299_/B _7048_/X _6947_/X _6943_/Y vssd1 vssd1 vccd1 vccd1 _7052_/B sky130_fd_sc_hd__o211ai_1
XFILLER_86_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6002_ _6002_/A _6221_/C vssd1 vssd1 vccd1 vccd1 _6004_/A sky130_fd_sc_hd__xnor2_1
XFILLER_94_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7953_ _8034_/A vssd1 vssd1 vccd1 vccd1 _8123_/S sky130_fd_sc_hd__buf_2
X_6904_ _6806_/A _6806_/B _6903_/X vssd1 vssd1 vccd1 vccd1 _6920_/A sky130_fd_sc_hd__a21o_1
XFILLER_82_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7884_ _7883_/B _7883_/C _7883_/A vssd1 vssd1 vccd1 vccd1 _7893_/B sky130_fd_sc_hd__a21o_1
XFILLER_23_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6835_ _6835_/A _6927_/A vssd1 vssd1 vccd1 vccd1 _6836_/B sky130_fd_sc_hd__nor2_2
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6766_ _6766_/A _6729_/A vssd1 vssd1 vccd1 vccd1 _6766_/X sky130_fd_sc_hd__or2b_1
XFILLER_50_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5717_ _5718_/A _5718_/B vssd1 vssd1 vccd1 vccd1 _5806_/B sky130_fd_sc_hd__nand2_1
X_8505_ _8505_/A _8505_/B vssd1 vssd1 vccd1 vccd1 _8505_/X sky130_fd_sc_hd__xor2_1
X_6697_ _6697_/A _6697_/B _6697_/C vssd1 vssd1 vccd1 vccd1 _6704_/A sky130_fd_sc_hd__nand3_1
XFILLER_40_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5648_ _5678_/A _5678_/B vssd1 vssd1 vccd1 vccd1 _5728_/A sky130_fd_sc_hd__and2b_1
X_8436_ _8429_/A _8434_/B _8429_/B vssd1 vssd1 vccd1 vccd1 _8493_/B sky130_fd_sc_hd__a21bo_1
X_8367_ _8367_/A vssd1 vssd1 vccd1 vccd1 _8367_/Y sky130_fd_sc_hd__inv_2
X_5579_ _6218_/A _5579_/B vssd1 vssd1 vccd1 vccd1 _5722_/A sky130_fd_sc_hd__xnor2_1
X_7318_ _7036_/A _7036_/B _7317_/Y vssd1 vssd1 vccd1 vccd1 _7319_/B sky130_fd_sc_hd__o21a_1
X_8298_ _8298_/A _8357_/B vssd1 vssd1 vccd1 vccd1 _8299_/B sky130_fd_sc_hd__xnor2_1
XFILLER_104_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7249_ _7249_/A _7286_/A vssd1 vssd1 vccd1 vccd1 _7289_/A sky130_fd_sc_hd__and2_1
XFILLER_104_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8789__56 vssd1 vssd1 vccd1 vccd1 _8789__56/HI _8898_/A sky130_fd_sc_hd__conb_1
XFILLER_92_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4950_ _5245_/A _4950_/B vssd1 vssd1 vccd1 vccd1 _5223_/D sky130_fd_sc_hd__nand2_2
X_4881_ _4957_/A _4891_/C _4990_/B vssd1 vssd1 vccd1 vccd1 _4890_/B sky130_fd_sc_hd__o21a_1
X_6620_ _6759_/A _6800_/A _6619_/Y vssd1 vssd1 vccd1 vccd1 _6916_/A sky130_fd_sc_hd__a21bo_1
X_6551_ _6590_/A vssd1 vssd1 vccd1 vccd1 _7065_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_20_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5502_ _5502_/A vssd1 vssd1 vccd1 vccd1 _5567_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6482_ _8714_/Q vssd1 vssd1 vccd1 vccd1 _7540_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5433_ _5427_/C _5432_/X _5433_/S vssd1 vssd1 vccd1 vccd1 _5434_/C sky130_fd_sc_hd__mux2_1
X_8221_ _8221_/A _8221_/B vssd1 vssd1 vccd1 vccd1 _8319_/B sky130_fd_sc_hd__xnor2_1
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8152_ _8152_/A _8152_/B vssd1 vssd1 vccd1 vccd1 _8155_/A sky130_fd_sc_hd__xor2_1
X_5364_ _8655_/Q vssd1 vssd1 vccd1 vccd1 _6353_/B sky130_fd_sc_hd__clkbuf_1
X_7103_ _7103_/A _7103_/B vssd1 vssd1 vccd1 vccd1 _7107_/A sky130_fd_sc_hd__or2_1
X_5295_ _8653_/Q _8652_/Q _5294_/X _8654_/Q vssd1 vssd1 vccd1 vccd1 _6502_/A sky130_fd_sc_hd__a31oi_1
X_8083_ _8108_/B _8083_/B vssd1 vssd1 vccd1 vccd1 _8096_/A sky130_fd_sc_hd__xnor2_1
X_7034_ _7034_/A _7034_/B vssd1 vssd1 vccd1 vccd1 _7317_/B sky130_fd_sc_hd__xnor2_1
XFILLER_87_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7936_ _7936_/A _7936_/B _7936_/C vssd1 vssd1 vccd1 vccd1 _7938_/A sky130_fd_sc_hd__nor3_1
X_7867_ _7867_/A _7867_/B _7867_/C vssd1 vssd1 vccd1 vccd1 _7881_/A sky130_fd_sc_hd__nand3_1
XFILLER_35_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6818_ _6818_/A _6818_/B vssd1 vssd1 vccd1 vccd1 _6819_/B sky130_fd_sc_hd__xor2_1
X_7798_ _8063_/A _7798_/B _7813_/B vssd1 vssd1 vccd1 vccd1 _7798_/X sky130_fd_sc_hd__and3_1
X_6749_ _7010_/A _7060_/B vssd1 vssd1 vccd1 vccd1 _7335_/B sky130_fd_sc_hd__nor2_4
XFILLER_7_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8419_ _8443_/A _8443_/B vssd1 vssd1 vccd1 vccd1 _8420_/B sky130_fd_sc_hd__xor2_2
XFILLER_2_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5080_ _5080_/A _5080_/B vssd1 vssd1 vccd1 vccd1 _5080_/Y sky130_fd_sc_hd__nor2_2
XFILLER_69_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5982_ _5983_/A _5983_/B vssd1 vssd1 vccd1 vccd1 _5982_/X sky130_fd_sc_hd__or2_1
X_4933_ _5245_/C vssd1 vssd1 vccd1 vccd1 _5044_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7721_ _7736_/A _8515_/B vssd1 vssd1 vccd1 vccd1 _7833_/A sky130_fd_sc_hd__nand2_1
XFILLER_32_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4864_ _4864_/A _4864_/B vssd1 vssd1 vccd1 vccd1 _4864_/X sky130_fd_sc_hd__and2_1
XFILLER_60_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7652_ _7652_/A _7652_/B vssd1 vssd1 vccd1 vccd1 _7741_/A sky130_fd_sc_hd__or2_1
X_6603_ _8713_/Q _6603_/B vssd1 vssd1 vccd1 vccd1 _6811_/B sky130_fd_sc_hd__nor2_1
X_4795_ _5591_/A _4795_/B _4795_/C vssd1 vssd1 vccd1 vccd1 _4796_/B sky130_fd_sc_hd__and3_1
XFILLER_20_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7583_ _8566_/S vssd1 vssd1 vccd1 vccd1 _8578_/A sky130_fd_sc_hd__clkbuf_2
X_6534_ _6534_/A _6541_/A vssd1 vssd1 vccd1 vccd1 _6538_/A sky130_fd_sc_hd__nand2_1
X_6465_ _6465_/A vssd1 vssd1 vccd1 vccd1 _8695_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5416_ _5415_/A _5415_/B _4581_/B vssd1 vssd1 vccd1 vccd1 _5416_/X sky130_fd_sc_hd__a21o_1
X_8204_ _8204_/A vssd1 vssd1 vccd1 vccd1 _8450_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6396_ _8694_/Q _6396_/B _8695_/Q _8693_/Q vssd1 vssd1 vccd1 vccd1 _6397_/C sky130_fd_sc_hd__and4b_1
X_5347_ _5351_/C _5347_/B vssd1 vssd1 vccd1 vccd1 _8648_/D sky130_fd_sc_hd__nor2_1
X_8135_ _8224_/A _8135_/B vssd1 vssd1 vccd1 vccd1 _8136_/B sky130_fd_sc_hd__nor2_1
XFILLER_87_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5278_ _8630_/Q _5285_/B vssd1 vssd1 vccd1 vccd1 _5278_/X sky130_fd_sc_hd__or2_1
X_8066_ _8066_/A _8146_/B vssd1 vssd1 vccd1 vccd1 _8370_/A sky130_fd_sc_hd__nand2_2
X_7017_ _7017_/A _7017_/B vssd1 vssd1 vccd1 vccd1 _7018_/C sky130_fd_sc_hd__xnor2_1
XFILLER_87_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8759__26 vssd1 vssd1 vccd1 vccd1 _8759__26/HI _8854_/A sky130_fd_sc_hd__conb_1
XFILLER_55_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7919_ _7919_/A _7919_/B vssd1 vssd1 vccd1 vccd1 _7920_/B sky130_fd_sc_hd__and2_1
XFILLER_102_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8899_ _8899_/A _4429_/Y vssd1 vssd1 vccd1 vccd1 io_out[36] sky130_fd_sc_hd__ebufn_8
XFILLER_62_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8773__40 vssd1 vssd1 vccd1 vccd1 _8773__40/HI _8868_/A sky130_fd_sc_hd__conb_1
XFILLER_61_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4580_ _5434_/B vssd1 vssd1 vccd1 vccd1 _4581_/B sky130_fd_sc_hd__clkbuf_2
X_6250_ _6250_/A _6250_/B vssd1 vssd1 vccd1 vccd1 _6251_/B sky130_fd_sc_hd__xnor2_1
X_5201_ _5103_/B _5199_/X _5200_/X _5143_/A vssd1 vssd1 vccd1 vccd1 _5205_/B sky130_fd_sc_hd__o211a_1
XFILLER_88_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6181_ _6181_/A _6181_/B vssd1 vssd1 vccd1 vccd1 _6182_/B sky130_fd_sc_hd__xor2_1
X_5132_ _5218_/A _5212_/B _5132_/C vssd1 vssd1 vccd1 vccd1 _5132_/X sky130_fd_sc_hd__or3_1
X_5063_ _5042_/X _5058_/X _5059_/X _5103_/A _4692_/A vssd1 vssd1 vccd1 vccd1 _5064_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_37_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5965_ _5906_/A _5965_/B vssd1 vssd1 vccd1 vccd1 _5965_/X sky130_fd_sc_hd__and2b_1
X_8684_ _8689_/CLK _8684_/D vssd1 vssd1 vccd1 vccd1 _8684_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4916_ _4916_/A _5188_/B _4991_/B _4916_/D vssd1 vssd1 vccd1 vccd1 _4916_/X sky130_fd_sc_hd__or4_1
X_5896_ _5896_/A _6001_/B vssd1 vssd1 vccd1 vccd1 _5899_/A sky130_fd_sc_hd__xnor2_1
X_7704_ _7712_/A _7712_/B vssd1 vssd1 vccd1 vccd1 _7859_/B sky130_fd_sc_hd__xor2_2
X_4847_ _4847_/A _4957_/A _4839_/B _4828_/A vssd1 vssd1 vccd1 vccd1 _4904_/A sky130_fd_sc_hd__or4bb_4
X_7635_ _7722_/A _7666_/B _7634_/X vssd1 vssd1 vccd1 vccd1 _7639_/A sky130_fd_sc_hd__a21o_1
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4778_ _4778_/A vssd1 vssd1 vccd1 vccd1 _8618_/D sky130_fd_sc_hd__clkbuf_1
X_7566_ _8571_/A _8576_/A _7564_/X _7565_/X _7499_/X vssd1 vssd1 vccd1 vccd1 _8716_/D
+ sky130_fd_sc_hd__o311ai_1
XFILLER_20_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6517_ _6509_/A _6526_/B _6510_/Y vssd1 vssd1 vccd1 vccd1 _6518_/B sky130_fd_sc_hd__a21o_1
X_7497_ _7491_/A _7491_/C _7491_/D _7496_/Y _7614_/A vssd1 vssd1 vccd1 vccd1 _7497_/X
+ sky130_fd_sc_hd__a41o_1
X_6448_ _6450_/B _6464_/B _6448_/C vssd1 vssd1 vccd1 vccd1 _6449_/A sky130_fd_sc_hd__and3b_1
X_6379_ _8685_/Q vssd1 vssd1 vccd1 vccd1 _6437_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8118_ _8118_/A _8118_/B _8118_/C vssd1 vssd1 vccd1 vccd1 _8131_/B sky130_fd_sc_hd__and3_1
XFILLER_102_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8049_ _8049_/A _8049_/B vssd1 vssd1 vccd1 vccd1 _8110_/B sky130_fd_sc_hd__xor2_2
XFILLER_90_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5750_ _5751_/A _5751_/C _5751_/B vssd1 vssd1 vccd1 vccd1 _5810_/A sky130_fd_sc_hd__a21oi_1
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4701_ _4697_/X _4700_/A _4700_/Y _4672_/X vssd1 vssd1 vccd1 vccd1 _8605_/D sky130_fd_sc_hd__o211a_1
X_5681_ _5967_/A vssd1 vssd1 vccd1 vccd1 _5943_/A sky130_fd_sc_hd__clkbuf_2
X_7420_ _7345_/A _7345_/B _7419_/X vssd1 vssd1 vccd1 vccd1 _7422_/A sky130_fd_sc_hd__a21oi_1
X_4632_ _8596_/Q _4632_/B vssd1 vssd1 vccd1 vccd1 _4637_/C sky130_fd_sc_hd__and2_1
X_7351_ _7351_/A _7351_/B vssd1 vssd1 vccd1 vccd1 _7364_/C sky130_fd_sc_hd__xnor2_1
X_4563_ _8627_/Q _4563_/B vssd1 vssd1 vccd1 vccd1 _4564_/A sky130_fd_sc_hd__and2_1
X_4494_ _7652_/B vssd1 vssd1 vccd1 vccd1 _4781_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7282_ _7495_/A _7493_/A _7493_/B _7278_/B _7278_/A vssd1 vssd1 vccd1 vccd1 _7469_/B
+ sky130_fd_sc_hd__o32a_1
X_6302_ _6302_/A _6302_/B vssd1 vssd1 vccd1 vccd1 _6320_/A sky130_fd_sc_hd__xor2_2
X_6233_ _6291_/A _6291_/B vssd1 vssd1 vccd1 vccd1 _6234_/B sky130_fd_sc_hd__xor2_4
XFILLER_69_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6164_ _5964_/A _5964_/B _6163_/X vssd1 vssd1 vccd1 vccd1 _6291_/A sky130_fd_sc_hd__a21oi_4
XFILLER_97_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5115_ _5115_/A _5192_/A _5188_/B _5227_/B vssd1 vssd1 vccd1 vccd1 _5237_/B sky130_fd_sc_hd__nor4_1
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6095_ _6095_/A vssd1 vssd1 vccd1 vccd1 _6095_/Y sky130_fd_sc_hd__clkinv_2
X_5046_ _5046_/A vssd1 vssd1 vccd1 vccd1 _5199_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6997_ _7364_/B _7443_/B vssd1 vssd1 vccd1 vccd1 _6997_/Y sky130_fd_sc_hd__nand2_1
X_5948_ _5948_/A _5948_/B vssd1 vssd1 vccd1 vccd1 _5952_/C sky130_fd_sc_hd__and2_1
XFILLER_43_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5879_ _5879_/A _5879_/B _5879_/C vssd1 vssd1 vccd1 vccd1 _5880_/B sky130_fd_sc_hd__or3_1
X_8667_ _8735_/CLK _8667_/D vssd1 vssd1 vccd1 vccd1 _8667_/Q sky130_fd_sc_hd__dfxtp_1
X_8598_ _8671_/CLK _8598_/D vssd1 vssd1 vccd1 vccd1 _8598_/Q sky130_fd_sc_hd__dfxtp_1
X_7618_ _7618_/A _7618_/B vssd1 vssd1 vccd1 vccd1 _7623_/B sky130_fd_sc_hd__or2_1
X_7549_ _7537_/C _7548_/C _7548_/A vssd1 vssd1 vccd1 vccd1 _7550_/C sky130_fd_sc_hd__o21ai_1
XFILLER_5_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_4_0_wb_clk_i clkbuf_4_5_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _8732_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_17_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8743__10 vssd1 vssd1 vccd1 vccd1 _8743__10/HI _8838_/A sky130_fd_sc_hd__conb_1
XFILLER_12_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6920_ _6920_/A _6920_/B vssd1 vssd1 vccd1 vccd1 _6921_/B sky130_fd_sc_hd__xor2_1
X_6851_ _7010_/A _7060_/B vssd1 vssd1 vccd1 vccd1 _7310_/A sky130_fd_sc_hd__or2_2
X_5802_ _5802_/A _5802_/B vssd1 vssd1 vccd1 vccd1 _5806_/A sky130_fd_sc_hd__or2_1
XFILLER_35_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6782_ _7350_/B vssd1 vssd1 vccd1 vccd1 _7352_/B sky130_fd_sc_hd__buf_2
XFILLER_50_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8521_ _8531_/A _8725_/Q vssd1 vssd1 vccd1 vccd1 _8521_/Y sky130_fd_sc_hd__nor2_1
X_5733_ _6120_/A _5833_/A _5962_/A vssd1 vssd1 vccd1 vccd1 _5841_/A sky130_fd_sc_hd__a21o_1
X_5664_ _5948_/B vssd1 vssd1 vccd1 vccd1 _6030_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_30_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8452_ _8452_/A _8452_/B vssd1 vssd1 vccd1 vccd1 _8453_/B sky130_fd_sc_hd__xnor2_1
X_7403_ _7403_/A _7403_/B vssd1 vssd1 vccd1 vccd1 _7405_/A sky130_fd_sc_hd__xnor2_1
X_4615_ _8590_/Q _4614_/B _4595_/X vssd1 vssd1 vccd1 vccd1 _4616_/B sky130_fd_sc_hd__o21ai_1
X_8383_ _8383_/A vssd1 vssd1 vccd1 vccd1 _8383_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5595_ _5595_/A _5595_/B vssd1 vssd1 vccd1 vccd1 _5948_/A sky130_fd_sc_hd__xnor2_4
X_7334_ _7434_/B _7454_/C vssd1 vssd1 vccd1 vccd1 _7338_/A sky130_fd_sc_hd__xor2_2
X_4546_ _8623_/Q _4552_/B vssd1 vssd1 vccd1 vccd1 _4547_/A sky130_fd_sc_hd__and2_1
X_7265_ _7270_/A _7270_/B _7264_/X vssd1 vssd1 vccd1 vccd1 _7286_/C sky130_fd_sc_hd__o21ai_1
XFILLER_1_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4477_ _7871_/A vssd1 vssd1 vccd1 vccd1 _6596_/B sky130_fd_sc_hd__clkbuf_4
X_7196_ _7430_/A _7409_/A _7196_/C vssd1 vssd1 vccd1 vccd1 _7196_/X sky130_fd_sc_hd__or3_1
X_6216_ _6005_/A _6005_/B _6215_/Y vssd1 vssd1 vccd1 vccd1 _6224_/A sky130_fd_sc_hd__a21o_1
XFILLER_85_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6147_ _6299_/A _6299_/C vssd1 vssd1 vccd1 vccd1 _6300_/B sky130_fd_sc_hd__or2_1
XFILLER_38_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_13 _8572_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6078_ _6111_/A vssd1 vssd1 vccd1 vccd1 _6078_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5029_ _5029_/A _5029_/B vssd1 vssd1 vccd1 vccd1 _5030_/A sky130_fd_sc_hd__or2_1
XFILLER_57_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8719_ _8735_/CLK _8719_/D vssd1 vssd1 vccd1 vccd1 _8719_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4400_ _4400_/A vssd1 vssd1 vccd1 vccd1 _4400_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5380_ _8662_/Q vssd1 vssd1 vccd1 vccd1 _5426_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4331_ input1/X vssd1 vssd1 vccd1 vccd1 _4456_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7050_ _6943_/Y _6947_/X _7048_/X _7299_/B vssd1 vssd1 vccd1 vccd1 _7050_/Y sky130_fd_sc_hd__a211oi_1
X_6001_ _6001_/A _6001_/B vssd1 vssd1 vccd1 vccd1 _6221_/C sky130_fd_sc_hd__xnor2_2
XFILLER_67_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7952_ _8139_/A _7952_/B vssd1 vssd1 vccd1 vccd1 _8034_/A sky130_fd_sc_hd__or2_1
X_6903_ _6816_/A _6903_/B vssd1 vssd1 vccd1 vccd1 _6903_/X sky130_fd_sc_hd__and2b_1
XFILLER_35_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7883_ _7883_/A _7883_/B _7883_/C vssd1 vssd1 vccd1 vccd1 _7893_/A sky130_fd_sc_hd__nand3_1
X_6834_ _6848_/A _6848_/B _6614_/A vssd1 vssd1 vccd1 vccd1 _6836_/A sky130_fd_sc_hd__a21o_2
XFILLER_62_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6765_ _6765_/A _6765_/B vssd1 vssd1 vccd1 vccd1 _7109_/B sky130_fd_sc_hd__xnor2_1
XFILLER_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5716_ _5716_/A _5802_/B vssd1 vssd1 vccd1 vccd1 _5718_/B sky130_fd_sc_hd__xnor2_1
X_8504_ _8506_/A _8506_/C _8506_/B vssd1 vssd1 vccd1 vccd1 _8505_/B sky130_fd_sc_hd__a21bo_1
X_6696_ _6804_/B _6696_/B vssd1 vssd1 vccd1 vccd1 _6697_/C sky130_fd_sc_hd__and2_1
X_8435_ _8496_/B _8496_/C _8497_/B _8496_/A vssd1 vssd1 vccd1 vccd1 _8493_/A sky130_fd_sc_hd__a211o_1
XFILLER_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5647_ _5685_/A _5687_/A vssd1 vssd1 vccd1 vccd1 _5678_/B sky130_fd_sc_hd__xnor2_1
X_8366_ _8066_/A _8072_/A _8166_/X _8365_/X vssd1 vssd1 vccd1 vccd1 _8372_/A sky130_fd_sc_hd__a31o_1
X_5578_ _5578_/A _5893_/B vssd1 vssd1 vccd1 vccd1 _5579_/B sky130_fd_sc_hd__xnor2_1
X_7317_ _7317_/A _7317_/B vssd1 vssd1 vccd1 vccd1 _7317_/Y sky130_fd_sc_hd__nand2_1
X_4529_ _7630_/B vssd1 vssd1 vccd1 vccd1 _4845_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_8297_ _8297_/A _8297_/B vssd1 vssd1 vccd1 vccd1 _8357_/B sky130_fd_sc_hd__xnor2_1
XFILLER_104_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7248_ _7249_/A _7248_/B _7248_/C vssd1 vssd1 vccd1 vccd1 _7286_/A sky130_fd_sc_hd__nand3_1
X_7179_ _7178_/A _7179_/B vssd1 vssd1 vccd1 vccd1 _7179_/X sky130_fd_sc_hd__and2b_1
XFILLER_58_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4880_ _5126_/A _5115_/A vssd1 vssd1 vccd1 vccd1 _5111_/A sky130_fd_sc_hd__or2_2
XFILLER_44_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6550_ _6593_/A _6593_/B vssd1 vssd1 vccd1 vccd1 _6590_/A sky130_fd_sc_hd__and2_1
XFILLER_20_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5501_ _5501_/A _5510_/C vssd1 vssd1 vccd1 vccd1 _6019_/A sky130_fd_sc_hd__xnor2_1
X_6481_ _8715_/Q _6481_/B _6500_/A vssd1 vssd1 vccd1 vccd1 _6481_/X sky130_fd_sc_hd__or3b_1
X_5432_ _5432_/A _5432_/B vssd1 vssd1 vccd1 vccd1 _5432_/X sky130_fd_sc_hd__or2_1
X_8220_ _8228_/A _8220_/B vssd1 vssd1 vccd1 vccd1 _8221_/B sky130_fd_sc_hd__xor2_1
X_5363_ _5361_/Y _5359_/C _5362_/X vssd1 vssd1 vccd1 vccd1 _8653_/D sky130_fd_sc_hd__a21boi_1
X_8151_ _8247_/B _8291_/A _8151_/S vssd1 vssd1 vccd1 vccd1 _8152_/B sky130_fd_sc_hd__mux2_1
XFILLER_99_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7102_ _7102_/A _7102_/B vssd1 vssd1 vccd1 vccd1 _7103_/B sky130_fd_sc_hd__and2_1
XFILLER_101_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5294_ _8651_/Q _8650_/Q _5294_/C vssd1 vssd1 vccd1 vccd1 _5294_/X sky130_fd_sc_hd__or3_1
X_8082_ _8082_/A _8082_/B vssd1 vssd1 vccd1 vccd1 _8083_/B sky130_fd_sc_hd__xnor2_1
XFILLER_101_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7033_ _7033_/A _7033_/B vssd1 vssd1 vccd1 vccd1 _7034_/B sky130_fd_sc_hd__xnor2_1
XFILLER_101_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7935_ _8015_/A _7935_/B vssd1 vssd1 vccd1 vccd1 _7936_/C sky130_fd_sc_hd__nand2_1
XFILLER_35_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7866_ _7887_/A _7887_/B _7865_/C _7865_/D vssd1 vssd1 vccd1 vccd1 _7867_/C sky130_fd_sc_hd__a22o_1
XFILLER_23_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6817_ _6924_/A _6924_/B vssd1 vssd1 vccd1 vccd1 _6818_/B sky130_fd_sc_hd__xor2_1
XFILLER_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7797_ _7851_/A _7851_/B vssd1 vssd1 vccd1 vccd1 _7825_/A sky130_fd_sc_hd__xnor2_1
X_6748_ _6748_/A _6748_/B vssd1 vssd1 vccd1 vccd1 _7060_/B sky130_fd_sc_hd__xnor2_4
X_6679_ _6722_/B vssd1 vssd1 vccd1 vccd1 _7169_/B sky130_fd_sc_hd__buf_2
X_8418_ _8418_/A _8418_/B vssd1 vssd1 vccd1 vccd1 _8443_/B sky130_fd_sc_hd__xnor2_1
X_8349_ _8383_/A _8349_/B vssd1 vssd1 vccd1 vccd1 _8359_/B sky130_fd_sc_hd__xnor2_1
XFILLER_104_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5981_ _5981_/A _5981_/B vssd1 vssd1 vccd1 vccd1 _5989_/A sky130_fd_sc_hd__nor2_1
XFILLER_37_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4932_ _4932_/A vssd1 vssd1 vccd1 vccd1 _5245_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_7720_ _8365_/A vssd1 vssd1 vccd1 vccd1 _8515_/B sky130_fd_sc_hd__clkbuf_2
X_7651_ _7652_/A _8619_/Q vssd1 vssd1 vccd1 vccd1 _7651_/X sky130_fd_sc_hd__and2_1
X_6602_ _8712_/Q _6746_/B vssd1 vssd1 vccd1 vccd1 _6602_/Y sky130_fd_sc_hd__nor2_1
X_4863_ _4863_/A vssd1 vssd1 vccd1 vccd1 _4920_/B sky130_fd_sc_hd__inv_2
X_4794_ _5591_/A _4822_/B vssd1 vssd1 vccd1 vccd1 _4823_/B sky130_fd_sc_hd__nor2_1
X_7582_ _8718_/Q vssd1 vssd1 vccd1 vccd1 _7630_/A sky130_fd_sc_hd__inv_2
X_6533_ _6536_/A vssd1 vssd1 vccd1 vccd1 _6533_/Y sky130_fd_sc_hd__inv_2
X_6464_ _6462_/Y _6464_/B vssd1 vssd1 vccd1 vccd1 _6465_/A sky130_fd_sc_hd__and2b_1
X_8203_ _8203_/A _8203_/B _8203_/C vssd1 vssd1 vccd1 vccd1 _8211_/A sky130_fd_sc_hd__and3_1
X_5415_ _5415_/A _5415_/B vssd1 vssd1 vccd1 vccd1 _5415_/Y sky130_fd_sc_hd__nor2_1
X_6395_ _6395_/A _6395_/B _6395_/C vssd1 vssd1 vccd1 vccd1 _6396_/B sky130_fd_sc_hd__and3_1
X_5346_ _8648_/Q _5344_/A _5323_/X vssd1 vssd1 vccd1 vccd1 _5347_/B sky130_fd_sc_hd__o21ai_1
X_8134_ _8224_/A _8135_/B vssd1 vssd1 vccd1 vccd1 _8211_/B sky130_fd_sc_hd__and2_2
XFILLER_99_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5277_ _8728_/Q _5271_/X _5276_/X _5267_/X vssd1 vssd1 vccd1 vccd1 _8629_/D sky130_fd_sc_hd__o211a_1
X_8065_ _8065_/A _8065_/B vssd1 vssd1 vccd1 vccd1 _8196_/A sky130_fd_sc_hd__nand2_2
X_7016_ _7306_/A _7016_/B vssd1 vssd1 vccd1 vccd1 _7017_/B sky130_fd_sc_hd__xnor2_1
XFILLER_83_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7918_ _7919_/A _7919_/B vssd1 vssd1 vccd1 vccd1 _8008_/B sky130_fd_sc_hd__nor2_1
XFILLER_43_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8898_ _8898_/A _4431_/Y vssd1 vssd1 vccd1 vccd1 io_out[35] sky130_fd_sc_hd__ebufn_8
XFILLER_70_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7849_ _7849_/A vssd1 vssd1 vccd1 vccd1 _8529_/A sky130_fd_sc_hd__inv_2
XFILLER_11_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5200_ _5200_/A _5200_/B _5200_/C _5229_/C vssd1 vssd1 vccd1 vccd1 _5200_/X sky130_fd_sc_hd__or4_1
X_6180_ _5958_/A _5958_/B _6179_/X vssd1 vssd1 vccd1 vccd1 _6181_/B sky130_fd_sc_hd__a21oi_1
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5131_ _5131_/A _5208_/C vssd1 vssd1 vccd1 vccd1 _5132_/C sky130_fd_sc_hd__or2_1
XFILLER_69_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5062_ _5106_/C _5154_/B _5062_/C vssd1 vssd1 vccd1 vccd1 _5103_/A sky130_fd_sc_hd__or3_1
XFILLER_57_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5964_ _5964_/A _5964_/B vssd1 vssd1 vccd1 vccd1 _6011_/A sky130_fd_sc_hd__xor2_1
X_7703_ _7711_/A _7703_/B vssd1 vssd1 vccd1 vccd1 _8515_/C sky130_fd_sc_hd__and2_1
X_8683_ _8689_/CLK _8683_/D vssd1 vssd1 vccd1 vccd1 _8683_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4915_ _5153_/A _5196_/B _5017_/C _5107_/C _4914_/X vssd1 vssd1 vccd1 vccd1 _4916_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_52_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5895_ _5713_/A _5885_/A _5569_/A vssd1 vssd1 vccd1 vccd1 _6001_/B sky130_fd_sc_hd__o21ba_2
XFILLER_33_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4846_ _4885_/B _4896_/A vssd1 vssd1 vccd1 vccd1 _5186_/C sky130_fd_sc_hd__nor2_1
X_7634_ _8719_/Q _8616_/Q vssd1 vssd1 vccd1 vccd1 _7634_/X sky130_fd_sc_hd__and2b_1
X_7565_ _7876_/A _7555_/A _8571_/B vssd1 vssd1 vccd1 vccd1 _7565_/X sky130_fd_sc_hd__a21bo_1
X_6516_ _6516_/A _6516_/B vssd1 vssd1 vccd1 vccd1 _6518_/A sky130_fd_sc_hd__nor2_1
X_4777_ _4781_/B _7537_/B _4777_/C vssd1 vssd1 vccd1 vccd1 _4778_/A sky130_fd_sc_hd__and3b_1
X_7496_ _7496_/A _7509_/A _7496_/C vssd1 vssd1 vccd1 vccd1 _7496_/Y sky130_fd_sc_hd__nor3_1
X_6447_ _6446_/B _8687_/Q _6441_/B _8689_/Q vssd1 vssd1 vccd1 vccd1 _6448_/C sky130_fd_sc_hd__a31o_1
X_6378_ _8690_/Q _8692_/Q _8691_/Q _8689_/Q vssd1 vssd1 vccd1 vccd1 _6395_/A sky130_fd_sc_hd__and4bb_1
X_8819__86 vssd1 vssd1 vccd1 vccd1 _8819__86/HI _8928_/A sky130_fd_sc_hd__conb_1
X_5329_ _6466_/D _5328_/C _8643_/Q vssd1 vssd1 vccd1 vccd1 _5330_/B sky130_fd_sc_hd__a21o_1
X_8117_ _8325_/A _8032_/B _8116_/X vssd1 vssd1 vccd1 vccd1 _8213_/A sky130_fd_sc_hd__a21bo_1
XFILLER_87_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8048_ _8139_/B _8045_/Y _8158_/A vssd1 vssd1 vccd1 vccd1 _8049_/B sky130_fd_sc_hd__a21oi_2
XFILLER_71_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4700_ _4700_/A _5056_/A vssd1 vssd1 vccd1 vccd1 _4700_/Y sky130_fd_sc_hd__nand2_1
X_5680_ _5680_/A _5680_/B vssd1 vssd1 vccd1 vccd1 _6026_/A sky130_fd_sc_hd__xnor2_1
X_4631_ _4631_/A vssd1 vssd1 vccd1 vccd1 _8595_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7350_ _7350_/A _7350_/B vssd1 vssd1 vccd1 vccd1 _7351_/B sky130_fd_sc_hd__xnor2_1
X_4562_ _4562_/A vssd1 vssd1 vccd1 vccd1 _8880_/A sky130_fd_sc_hd__clkbuf_1
X_7281_ _6592_/A _6592_/B _7280_/X vssd1 vssd1 vccd1 vccd1 _7493_/B sky130_fd_sc_hd__a21oi_2
X_4493_ _8619_/Q vssd1 vssd1 vccd1 vccd1 _7652_/B sky130_fd_sc_hd__buf_2
X_6301_ _6296_/X _6332_/A _6300_/X vssd1 vssd1 vccd1 vccd1 _6315_/A sky130_fd_sc_hd__o21a_1
X_6232_ _6232_/A _6232_/B vssd1 vssd1 vccd1 vccd1 _6291_/B sky130_fd_sc_hd__xnor2_2
XFILLER_97_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6163_ _5963_/A _6163_/B vssd1 vssd1 vccd1 vccd1 _6163_/X sky130_fd_sc_hd__and2b_1
XFILLER_84_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5114_ _5114_/A vssd1 vssd1 vccd1 vccd1 _5227_/B sky130_fd_sc_hd__clkbuf_2
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6094_ _6094_/A _6094_/B vssd1 vssd1 vccd1 vccd1 _6306_/A sky130_fd_sc_hd__nor2_1
X_5045_ _5154_/B _5045_/B vssd1 vssd1 vccd1 vccd1 _5045_/X sky130_fd_sc_hd__or2_1
XFILLER_84_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6996_ _6918_/A _6918_/B _6995_/X vssd1 vssd1 vccd1 vccd1 _7017_/A sky130_fd_sc_hd__o21ai_1
XFILLER_80_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5947_ _5948_/A _5948_/B vssd1 vssd1 vccd1 vccd1 _5947_/X sky130_fd_sc_hd__or2_1
XFILLER_43_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8735_ _8735_/CLK _8735_/D vssd1 vssd1 vccd1 vccd1 _8735_/Q sky130_fd_sc_hd__dfxtp_1
X_8666_ _8732_/CLK _8666_/D vssd1 vssd1 vccd1 vccd1 _8666_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5878_ _5879_/A _5879_/B _5879_/C vssd1 vssd1 vccd1 vccd1 _5978_/A sky130_fd_sc_hd__o21ai_2
XFILLER_21_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7617_ _7618_/A _7617_/B vssd1 vssd1 vccd1 vccd1 _7619_/A sky130_fd_sc_hd__nand2_1
X_4829_ _4879_/B _4849_/B vssd1 vssd1 vccd1 vccd1 _5244_/B sky130_fd_sc_hd__nor2_2
X_8597_ _8600_/CLK _8597_/D vssd1 vssd1 vccd1 vccd1 _8597_/Q sky130_fd_sc_hd__dfxtp_1
X_7548_ _7548_/A _7548_/B _7548_/C vssd1 vssd1 vccd1 vccd1 _7550_/B sky130_fd_sc_hd__or3_1
X_7479_ _7479_/A _7479_/B vssd1 vssd1 vccd1 vccd1 _7480_/B sky130_fd_sc_hd__nand2_1
XFILLER_68_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6850_ _6929_/B vssd1 vssd1 vccd1 vccd1 _6926_/A sky130_fd_sc_hd__buf_2
XFILLER_35_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6781_ _7169_/B _7083_/B _6716_/X _6725_/B _6780_/Y vssd1 vssd1 vccd1 vccd1 _6905_/A
+ sky130_fd_sc_hd__a32oi_4
XFILLER_50_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5801_ _5801_/A _5870_/B vssd1 vssd1 vccd1 vccd1 _5808_/A sky130_fd_sc_hd__xnor2_1
X_5732_ _5732_/A _5742_/A vssd1 vssd1 vccd1 vccd1 _6273_/S sky130_fd_sc_hd__nand2_1
X_8520_ _8525_/B _8520_/B _7846_/Y vssd1 vssd1 vccd1 vccd1 _8520_/X sky130_fd_sc_hd__or3b_2
X_5663_ _5663_/A _5663_/B vssd1 vssd1 vccd1 vccd1 _5948_/B sky130_fd_sc_hd__or2_1
X_8451_ _8450_/B _8450_/C _8450_/Y vssd1 vssd1 vccd1 vccd1 _8452_/B sky130_fd_sc_hd__a21oi_1
X_7402_ _7403_/A _7320_/B _7401_/X vssd1 vssd1 vccd1 vccd1 _7403_/B sky130_fd_sc_hd__a21o_1
X_4614_ _8590_/Q _4614_/B vssd1 vssd1 vccd1 vccd1 _4619_/C sky130_fd_sc_hd__and2_1
X_8382_ _8382_/A _8382_/B vssd1 vssd1 vccd1 vccd1 _8423_/A sky130_fd_sc_hd__xnor2_1
X_5594_ _5594_/A _5594_/B vssd1 vssd1 vccd1 vccd1 _5595_/B sky130_fd_sc_hd__nor2_2
X_4545_ _4545_/A vssd1 vssd1 vccd1 vccd1 _8876_/A sky130_fd_sc_hd__clkbuf_1
X_7333_ _7333_/A vssd1 vssd1 vccd1 vccd1 _7454_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_104_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7264_ _7264_/A _7264_/B vssd1 vssd1 vccd1 vccd1 _7264_/X sky130_fd_sc_hd__or2_1
X_4476_ _8611_/Q vssd1 vssd1 vccd1 vccd1 _7871_/A sky130_fd_sc_hd__buf_2
X_7195_ _7195_/A _7195_/B vssd1 vssd1 vccd1 vccd1 _7198_/B sky130_fd_sc_hd__xnor2_1
X_6215_ _6215_/A _6215_/B vssd1 vssd1 vccd1 vccd1 _6215_/Y sky130_fd_sc_hd__nor2_1
X_6146_ _6146_/A _6146_/B vssd1 vssd1 vccd1 vccd1 _6299_/A sky130_fd_sc_hd__nand2_1
XFILLER_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_14 _8576_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6077_ _6110_/A _6110_/B vssd1 vssd1 vccd1 vccd1 _6111_/A sky130_fd_sc_hd__nor2_1
XFILLER_85_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5028_ _5190_/A _5028_/B _5028_/C vssd1 vssd1 vccd1 vccd1 _5028_/X sky130_fd_sc_hd__or3_1
XFILLER_72_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6979_ _6978_/A _6978_/B _6978_/C vssd1 vssd1 vccd1 vccd1 _6985_/B sky130_fd_sc_hd__a21o_1
X_8718_ _8732_/CLK _8718_/D vssd1 vssd1 vccd1 vccd1 _8718_/Q sky130_fd_sc_hd__dfxtp_1
X_8649_ _8677_/CLK _8649_/D vssd1 vssd1 vccd1 vccd1 _8649_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8803__70 vssd1 vssd1 vccd1 vccd1 _8803__70/HI _8912_/A sky130_fd_sc_hd__conb_1
XFILLER_17_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6000_ _6000_/A _6000_/B vssd1 vssd1 vccd1 vccd1 _6005_/A sky130_fd_sc_hd__xor2_2
XFILLER_67_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7951_ _7886_/A _7887_/B _7865_/C _7950_/X vssd1 vssd1 vccd1 vccd1 _7958_/A sky130_fd_sc_hd__a31o_1
XFILLER_27_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6902_ _6902_/A _6902_/B vssd1 vssd1 vccd1 vccd1 _6950_/A sky130_fd_sc_hd__nand2_1
X_7882_ _7881_/A _7881_/B _7881_/C vssd1 vssd1 vccd1 vccd1 _7883_/C sky130_fd_sc_hd__a21o_1
XFILLER_54_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6833_ _6857_/A _6857_/B vssd1 vssd1 vccd1 vccd1 _6833_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_23_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6764_ _7099_/B _6845_/B vssd1 vssd1 vccd1 vccd1 _6765_/B sky130_fd_sc_hd__xnor2_1
X_6695_ _6694_/B _6672_/A _6724_/A vssd1 vssd1 vccd1 vccd1 _6696_/B sky130_fd_sc_hd__a21o_1
XFILLER_50_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5715_ _5571_/A _5571_/B _5569_/X vssd1 vssd1 vccd1 vccd1 _5802_/B sky130_fd_sc_hd__a21oi_1
X_8503_ _8503_/A _8503_/B vssd1 vssd1 vccd1 vccd1 _8505_/A sky130_fd_sc_hd__xnor2_1
X_5646_ _5962_/A _5640_/Y _6049_/A vssd1 vssd1 vccd1 vccd1 _5687_/A sky130_fd_sc_hd__a21oi_2
X_8434_ _8497_/A _8434_/B vssd1 vssd1 vccd1 vccd1 _8496_/A sky130_fd_sc_hd__nand2_1
X_8365_ _8365_/A _8365_/B _8365_/C vssd1 vssd1 vccd1 vccd1 _8365_/X sky130_fd_sc_hd__and3_1
X_5577_ _5531_/A _6218_/A _5532_/B _5532_/A vssd1 vssd1 vccd1 vccd1 _5580_/A sky130_fd_sc_hd__a22o_1
X_7316_ _7316_/A _7316_/B vssd1 vssd1 vccd1 vccd1 _7401_/B sky130_fd_sc_hd__xor2_1
X_4528_ _6596_/B _6605_/B vssd1 vssd1 vccd1 vccd1 _4668_/A sky130_fd_sc_hd__nand2_1
X_8296_ _8296_/A _8296_/B vssd1 vssd1 vccd1 vccd1 _8297_/B sky130_fd_sc_hd__nor2_1
X_4459_ _4461_/A vssd1 vssd1 vccd1 vccd1 _4459_/Y sky130_fd_sc_hd__inv_2
X_7247_ _7245_/A _7245_/C _7245_/B vssd1 vssd1 vccd1 vccd1 _7248_/C sky130_fd_sc_hd__a21o_1
XFILLER_49_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7178_ _7178_/A _7179_/B vssd1 vssd1 vccd1 vccd1 _7187_/B sky130_fd_sc_hd__xnor2_1
XFILLER_85_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6129_ _6129_/A _6129_/B vssd1 vssd1 vccd1 vccd1 _6130_/B sky130_fd_sc_hd__and2_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5500_ _5500_/A _5500_/B vssd1 vssd1 vccd1 vccd1 _5510_/C sky130_fd_sc_hd__xor2_1
X_6480_ _7520_/A _7514_/A _7526_/A vssd1 vssd1 vccd1 vccd1 _6481_/B sky130_fd_sc_hd__o21a_1
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5431_ _8663_/Q vssd1 vssd1 vccd1 vccd1 _5634_/A sky130_fd_sc_hd__clkinv_2
X_5362_ _5362_/A vssd1 vssd1 vccd1 vccd1 _5362_/X sky130_fd_sc_hd__buf_2
X_8150_ _8150_/A _8304_/A vssd1 vssd1 vccd1 vccd1 _8151_/S sky130_fd_sc_hd__nor2_1
XFILLER_99_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7101_ _7101_/A _7101_/B vssd1 vssd1 vccd1 vccd1 _7127_/B sky130_fd_sc_hd__xnor2_2
X_8081_ _8081_/A _8081_/B vssd1 vssd1 vccd1 vccd1 _8082_/B sky130_fd_sc_hd__xnor2_2
X_5293_ _8647_/Q _5292_/X _8649_/Q _8648_/Q vssd1 vssd1 vccd1 vccd1 _5294_/C sky130_fd_sc_hd__o211a_1
X_7032_ _7335_/B _7032_/B vssd1 vssd1 vccd1 vccd1 _7033_/B sky130_fd_sc_hd__xnor2_1
XFILLER_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7934_ _7934_/A _7934_/B vssd1 vssd1 vccd1 vccd1 _7935_/B sky130_fd_sc_hd__nand2_1
X_8794__61 vssd1 vssd1 vccd1 vccd1 _8794__61/HI _8903_/A sky130_fd_sc_hd__conb_1
XFILLER_82_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7865_ _7886_/A _7887_/B _7865_/C _7865_/D vssd1 vssd1 vccd1 vccd1 _7867_/B sky130_fd_sc_hd__nand4_1
XFILLER_51_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6816_ _6816_/A _6903_/B vssd1 vssd1 vccd1 vccd1 _6924_/B sky130_fd_sc_hd__xor2_1
X_7796_ _8399_/A _8515_/D _7796_/C vssd1 vssd1 vccd1 vccd1 _7851_/B sky130_fd_sc_hd__or3_1
X_6747_ _6747_/A _6747_/B vssd1 vssd1 vccd1 vccd1 _6748_/B sky130_fd_sc_hd__nand2_2
XFILLER_11_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6678_ _6678_/A _6678_/B vssd1 vssd1 vccd1 vccd1 _6722_/B sky130_fd_sc_hd__xor2_1
X_5629_ _5682_/A _5676_/B _5628_/X vssd1 vssd1 vccd1 vccd1 _5678_/A sky130_fd_sc_hd__a21oi_1
X_8417_ _8414_/A _8414_/B _8416_/X vssd1 vssd1 vccd1 vccd1 _8418_/B sky130_fd_sc_hd__a21oi_1
X_8348_ _8384_/A _8384_/B vssd1 vssd1 vccd1 vccd1 _8349_/B sky130_fd_sc_hd__xor2_1
XFILLER_2_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8279_ _8489_/A _8279_/B vssd1 vssd1 vccd1 vccd1 _8279_/Y sky130_fd_sc_hd__nor2_1
XFILLER_76_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5980_ _5978_/A _5880_/B _5905_/B _5904_/B _5904_/A vssd1 vssd1 vccd1 vccd1 _6188_/A
+ sky130_fd_sc_hd__a32o_1
X_4931_ _5200_/A vssd1 vssd1 vccd1 vccd1 _5171_/C sky130_fd_sc_hd__clkbuf_2
X_4862_ _4868_/A vssd1 vssd1 vccd1 vccd1 _4903_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_17_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7650_ _7642_/A _7642_/B _7644_/X _7645_/A vssd1 vssd1 vccd1 vccd1 _7654_/A sky130_fd_sc_hd__a31o_1
X_6601_ _6593_/A _6582_/B _6558_/B _6553_/X vssd1 vssd1 vccd1 vccd1 _6745_/B sky130_fd_sc_hd__a211o_1
XFILLER_60_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4793_ _4822_/A _4822_/B vssd1 vssd1 vccd1 vccd1 _4859_/A sky130_fd_sc_hd__nor2_1
X_7581_ _7617_/B _7555_/Y _7578_/Y _7580_/X _7544_/X vssd1 vssd1 vccd1 vccd1 _8717_/D
+ sky130_fd_sc_hd__a221o_1
X_6532_ _6508_/A _6541_/A _6529_/X _6531_/X vssd1 vssd1 vccd1 vccd1 _8702_/D sky130_fd_sc_hd__a31o_1
X_6463_ _8694_/Q _6461_/A _6462_/Y _4746_/X vssd1 vssd1 vccd1 vccd1 _8694_/D sky130_fd_sc_hd__o211a_1
X_8202_ _8143_/A _8143_/B _8201_/X vssd1 vssd1 vccd1 vccd1 _8239_/A sky130_fd_sc_hd__a21oi_1
X_5414_ _5406_/B _5408_/B _5406_/A vssd1 vssd1 vccd1 vccd1 _5415_/B sky130_fd_sc_hd__o21ba_1
X_6394_ _8680_/Q _8686_/Q _8685_/Q _6394_/D vssd1 vssd1 vccd1 vccd1 _6395_/C sky130_fd_sc_hd__and4bb_1
X_8133_ _8133_/A _8203_/C vssd1 vssd1 vccd1 vccd1 _8135_/B sky130_fd_sc_hd__xnor2_1
X_5345_ _8648_/Q _8647_/Q _5345_/C vssd1 vssd1 vccd1 vccd1 _5351_/C sky130_fd_sc_hd__and3_1
XFILLER_101_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5276_ _8629_/Q _5276_/B vssd1 vssd1 vccd1 vccd1 _5276_/X sky130_fd_sc_hd__or2_1
X_8064_ _8309_/A vssd1 vssd1 vccd1 vccd1 _8291_/A sky130_fd_sc_hd__clkbuf_2
X_7015_ _7015_/A _7015_/B vssd1 vssd1 vccd1 vccd1 _7016_/B sky130_fd_sc_hd__xnor2_1
XFILLER_87_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7917_ _7903_/C _7814_/B _7649_/B _8308_/A vssd1 vssd1 vccd1 vccd1 _7919_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_43_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8897_ _8897_/A _4463_/Y vssd1 vssd1 vccd1 vccd1 io_out[34] sky130_fd_sc_hd__ebufn_8
XFILLER_70_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7848_ _7848_/A _7848_/B vssd1 vssd1 vccd1 vccd1 _7849_/A sky130_fd_sc_hd__and2_1
X_7779_ _7779_/A _7886_/C vssd1 vssd1 vccd1 vccd1 _7780_/B sky130_fd_sc_hd__xnor2_1
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5130_ _5130_/A _5171_/C vssd1 vssd1 vccd1 vccd1 _5218_/D sky130_fd_sc_hd__or2_1
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5061_ _5231_/B vssd1 vssd1 vccd1 vccd1 _5106_/C sky130_fd_sc_hd__buf_2
XFILLER_84_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5963_ _5963_/A _6163_/B vssd1 vssd1 vccd1 vccd1 _5964_/B sky130_fd_sc_hd__xnor2_2
XFILLER_25_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8764__31 vssd1 vssd1 vccd1 vccd1 _8764__31/HI _8859_/A sky130_fd_sc_hd__conb_1
X_4914_ _4914_/A _5115_/A vssd1 vssd1 vccd1 vccd1 _4914_/X sky130_fd_sc_hd__or2_1
XFILLER_18_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7702_ _7886_/A vssd1 vssd1 vccd1 vccd1 _8515_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_8682_ _8689_/CLK _8682_/D vssd1 vssd1 vccd1 vccd1 _8682_/Q sky130_fd_sc_hd__dfxtp_1
X_5894_ _5798_/A _6211_/B _5790_/A _6221_/A vssd1 vssd1 vccd1 vccd1 _5901_/B sky130_fd_sc_hd__o211a_1
X_4845_ _4845_/A _4845_/B _4845_/C _8612_/Q vssd1 vssd1 vccd1 vccd1 _4896_/A sky130_fd_sc_hd__or4_4
X_7633_ _8719_/Q _8616_/Q vssd1 vssd1 vccd1 vccd1 _7666_/B sky130_fd_sc_hd__xnor2_4
X_4776_ _4774_/B _4774_/C _4799_/A vssd1 vssd1 vccd1 vccd1 _4777_/C sky130_fd_sc_hd__a21o_1
X_7564_ _7876_/A _7555_/Y _7557_/X _7563_/X vssd1 vssd1 vccd1 vccd1 _7564_/X sky130_fd_sc_hd__o31a_1
X_6515_ _6515_/A _6515_/B vssd1 vssd1 vccd1 vccd1 _6516_/B sky130_fd_sc_hd__and2_1
X_7495_ _7495_/A _7501_/B vssd1 vssd1 vccd1 vccd1 _7496_/C sky130_fd_sc_hd__nor2_1
X_6446_ _8689_/Q _6446_/B _6446_/C vssd1 vssd1 vccd1 vccd1 _6450_/B sky130_fd_sc_hd__and3_1
X_6377_ _8691_/Q vssd1 vssd1 vccd1 vccd1 _6455_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_102_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5328_ _8643_/Q _8642_/Q _5328_/C vssd1 vssd1 vccd1 vccd1 _5332_/B sky130_fd_sc_hd__and3_1
X_8116_ _8116_/A _8031_/A vssd1 vssd1 vccd1 vccd1 _8116_/X sky130_fd_sc_hd__or2b_1
XFILLER_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8047_ _8045_/Y _8046_/X _8139_/B vssd1 vssd1 vccd1 vccd1 _8158_/A sky130_fd_sc_hd__a21oi_2
XFILLER_102_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5259_ _8622_/Q _5263_/B vssd1 vssd1 vccd1 vccd1 _5259_/X sky130_fd_sc_hd__or2_1
XFILLER_87_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4630_ _4632_/B _4645_/B _4630_/C vssd1 vssd1 vccd1 vccd1 _4631_/A sky130_fd_sc_hd__and3b_1
XFILLER_30_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4561_ _8626_/Q _4563_/B vssd1 vssd1 vccd1 vccd1 _4562_/A sky130_fd_sc_hd__and2_1
XFILLER_8_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6300_ _6311_/A _6300_/B _6300_/C vssd1 vssd1 vccd1 vccd1 _6300_/X sky130_fd_sc_hd__and3b_1
X_7280_ _7280_/A _7280_/B _7280_/C vssd1 vssd1 vccd1 vccd1 _7280_/X sky130_fd_sc_hd__and3_1
X_4492_ _4795_/B vssd1 vssd1 vccd1 vccd1 _4765_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6231_ _6231_/A _6283_/B vssd1 vssd1 vccd1 vccd1 _6232_/B sky130_fd_sc_hd__xnor2_4
XFILLER_103_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6162_ _6013_/A _6013_/B _6161_/X vssd1 vssd1 vccd1 vccd1 _6234_/A sky130_fd_sc_hd__a21o_2
XFILLER_97_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5113_ _4923_/X _5218_/A _5202_/D _5136_/C _5112_/X vssd1 vssd1 vccd1 vccd1 _5113_/X
+ sky130_fd_sc_hd__o32a_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6093_ _6157_/A _6092_/B _6090_/X vssd1 vssd1 vccd1 vccd1 _6094_/B sky130_fd_sc_hd__a21boi_1
X_5044_ _5120_/A _5044_/B _5044_/C _5143_/B vssd1 vssd1 vccd1 vccd1 _5045_/B sky130_fd_sc_hd__or4_1
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6995_ _6995_/A _6995_/B vssd1 vssd1 vccd1 vccd1 _6995_/X sky130_fd_sc_hd__or2_1
XFILLER_53_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8734_ _8734_/CLK _8734_/D vssd1 vssd1 vccd1 vccd1 _8734_/Q sky130_fd_sc_hd__dfxtp_1
X_5946_ _5863_/B _5973_/A _5956_/B _5970_/B vssd1 vssd1 vccd1 vccd1 _6168_/A sky130_fd_sc_hd__a22oi_4
XFILLER_25_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5877_ _5981_/A _6265_/A _5981_/B vssd1 vssd1 vccd1 vccd1 _5879_/C sky130_fd_sc_hd__mux2_1
X_8665_ _8732_/CLK _8665_/D vssd1 vssd1 vccd1 vccd1 _8665_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4828_ _4828_/A _4847_/A _4828_/C vssd1 vssd1 vccd1 vccd1 _4879_/B sky130_fd_sc_hd__or3_2
X_7616_ _7613_/A _7613_/C _7613_/B vssd1 vssd1 vccd1 vccd1 _7620_/A sky130_fd_sc_hd__a21bo_1
X_8596_ _8600_/CLK _8596_/D vssd1 vssd1 vccd1 vccd1 _8596_/Q sky130_fd_sc_hd__dfxtp_1
X_7547_ _7539_/Y _7546_/X _7547_/S vssd1 vssd1 vccd1 vccd1 _7548_/C sky130_fd_sc_hd__mux2_1
X_4759_ _4758_/A _4758_/B _4752_/X vssd1 vssd1 vccd1 vccd1 _4759_/X sky130_fd_sc_hd__o21ba_1
X_7478_ _7478_/A _7482_/A vssd1 vssd1 vccd1 vccd1 _7480_/A sky130_fd_sc_hd__nand2_1
XFILLER_4_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6429_ _8683_/Q _6432_/C vssd1 vssd1 vccd1 vccd1 _6431_/A sky130_fd_sc_hd__and2_1
XFILLER_68_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6780_ _6780_/A _6780_/B vssd1 vssd1 vccd1 vccd1 _6780_/Y sky130_fd_sc_hd__nand2_1
X_5800_ _5800_/A _5800_/B vssd1 vssd1 vccd1 vccd1 _5870_/B sky130_fd_sc_hd__xnor2_1
XFILLER_62_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5731_ _6030_/A _6097_/B vssd1 vssd1 vccd1 vccd1 _5941_/B sky130_fd_sc_hd__nand2_1
X_5662_ _5661_/A _5661_/B _5661_/C vssd1 vssd1 vccd1 vccd1 _5663_/B sky130_fd_sc_hd__a21oi_2
X_8450_ _8450_/A _8450_/B _8450_/C vssd1 vssd1 vccd1 vccd1 _8450_/Y sky130_fd_sc_hd__nor3_1
X_7401_ _7319_/B _7401_/B vssd1 vssd1 vccd1 vccd1 _7401_/X sky130_fd_sc_hd__and2b_1
X_8381_ _8381_/A vssd1 vssd1 vccd1 vccd1 _8382_/B sky130_fd_sc_hd__inv_2
X_5593_ _8659_/Q _8617_/Q vssd1 vssd1 vccd1 vccd1 _5594_/B sky130_fd_sc_hd__and2b_1
X_4613_ _4613_/A vssd1 vssd1 vccd1 vccd1 _8589_/D sky130_fd_sc_hd__clkbuf_1
X_7332_ _7332_/A _7332_/B vssd1 vssd1 vccd1 vccd1 _7333_/A sky130_fd_sc_hd__or2_1
X_4544_ _8622_/Q _4552_/B vssd1 vssd1 vccd1 vccd1 _4545_/A sky130_fd_sc_hd__and2_2
X_7263_ _7264_/A _7264_/B vssd1 vssd1 vccd1 vccd1 _7270_/B sky130_fd_sc_hd__xnor2_2
XFILLER_104_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4475_ _4480_/C _4662_/A vssd1 vssd1 vccd1 vccd1 _4479_/C sky130_fd_sc_hd__nor2_1
X_6214_ _6221_/B _6221_/C vssd1 vssd1 vccd1 vccd1 _6215_/A sky130_fd_sc_hd__xnor2_1
X_7194_ _7225_/A _7225_/B _7193_/A vssd1 vssd1 vccd1 vccd1 _7198_/A sky130_fd_sc_hd__o21bai_1
X_6145_ _6299_/B _6299_/C vssd1 vssd1 vccd1 vccd1 _6311_/A sky130_fd_sc_hd__nor2_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_15 _7614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6076_ _6082_/A _6076_/B vssd1 vssd1 vccd1 vccd1 _6110_/B sky130_fd_sc_hd__nand2_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5027_ _5106_/B _5230_/B _5027_/C vssd1 vssd1 vccd1 vccd1 _5028_/C sky130_fd_sc_hd__or3_1
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6978_ _6978_/A _6978_/B _6978_/C vssd1 vssd1 vccd1 vccd1 _6985_/A sky130_fd_sc_hd__nand3_1
X_8717_ _8732_/CLK _8717_/D vssd1 vssd1 vccd1 vccd1 _8717_/Q sky130_fd_sc_hd__dfxtp_1
X_5929_ _6060_/A _6060_/B _6060_/C vssd1 vssd1 vccd1 vccd1 _6061_/A sky130_fd_sc_hd__o21a_1
XFILLER_41_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8648_ _8677_/CLK _8648_/D vssd1 vssd1 vccd1 vccd1 _8648_/Q sky130_fd_sc_hd__dfxtp_1
X_8579_ _7876_/A _8578_/Y _8531_/A vssd1 vssd1 vccd1 vccd1 _8579_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7950_ _7950_/A _7950_/B vssd1 vssd1 vccd1 vccd1 _7950_/X sky130_fd_sc_hd__and2_1
XFILLER_94_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6901_ _6901_/A _6901_/B _6901_/C vssd1 vssd1 vccd1 vccd1 _6902_/B sky130_fd_sc_hd__nand3_1
X_7881_ _7881_/A _7881_/B _7881_/C vssd1 vssd1 vccd1 vccd1 _7883_/B sky130_fd_sc_hd__nand3_1
X_6832_ _7196_/C _6839_/B _6831_/Y vssd1 vssd1 vccd1 vccd1 _6857_/B sky130_fd_sc_hd__a21oi_1
XFILLER_62_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6763_ _6763_/A _6763_/B vssd1 vssd1 vccd1 vccd1 _6845_/B sky130_fd_sc_hd__xnor2_1
XFILLER_50_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6694_ _6724_/A _6694_/B _6804_/A vssd1 vssd1 vccd1 vccd1 _6804_/B sky130_fd_sc_hd__nand3_1
X_5714_ _5578_/A _5788_/B _5579_/B _5713_/X vssd1 vssd1 vccd1 vccd1 _5718_/A sky130_fd_sc_hd__a22o_1
X_8502_ _8501_/B _8510_/A _8501_/A vssd1 vssd1 vccd1 vccd1 _8502_/Y sky130_fd_sc_hd__o21ai_1
X_5645_ _5641_/Y _5614_/B _5859_/A _5910_/B vssd1 vssd1 vccd1 vccd1 _6049_/A sky130_fd_sc_hd__o211a_1
X_8433_ _8433_/A _8433_/B vssd1 vssd1 vccd1 vccd1 _8434_/B sky130_fd_sc_hd__or2_1
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8364_ _8314_/A _8314_/B _8312_/Y vssd1 vssd1 vccd1 vccd1 _8373_/A sky130_fd_sc_hd__a21oi_1
X_5576_ _5713_/A vssd1 vssd1 vccd1 vccd1 _6218_/A sky130_fd_sc_hd__buf_2
X_7315_ _7315_/A _7315_/B vssd1 vssd1 vccd1 vccd1 _7316_/B sky130_fd_sc_hd__nand2_1
X_4527_ _4480_/C _4524_/X _4662_/A _4733_/S _4801_/B vssd1 vssd1 vccd1 vccd1 _4527_/X
+ sky130_fd_sc_hd__a2111o_1
X_8295_ _8295_/A _8295_/B _8295_/C vssd1 vssd1 vccd1 vccd1 _8296_/B sky130_fd_sc_hd__and3_1
XFILLER_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4458_ _4461_/A vssd1 vssd1 vccd1 vccd1 _4458_/Y sky130_fd_sc_hd__inv_2
X_7246_ _7010_/B _6926_/A _7165_/B _7173_/A vssd1 vssd1 vccd1 vccd1 _7248_/B sky130_fd_sc_hd__a2bb2o_1
X_7177_ _7177_/A _7177_/B vssd1 vssd1 vccd1 vccd1 _7179_/B sky130_fd_sc_hd__xor2_1
XFILLER_98_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4389_ _4401_/A vssd1 vssd1 vccd1 vccd1 _4394_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_58_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6128_ _6129_/A _6129_/B vssd1 vssd1 vccd1 vccd1 _6130_/A sky130_fd_sc_hd__nor2_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6059_ _6091_/A _6091_/B _6091_/C vssd1 vssd1 vccd1 vccd1 _6157_/A sky130_fd_sc_hd__o21ai_2
XFILLER_45_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5430_ _5398_/X _5429_/X _5426_/A _4582_/B vssd1 vssd1 vccd1 vccd1 _8662_/D sky130_fd_sc_hd__o2bb2a_1
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5361_ _8653_/Q vssd1 vssd1 vccd1 vccd1 _5361_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5292_ _8645_/Q _8644_/Q _5291_/X _8646_/Q vssd1 vssd1 vccd1 vccd1 _5292_/X sky130_fd_sc_hd__a31o_1
X_7100_ _7099_/B _7099_/C _7099_/A vssd1 vssd1 vccd1 vccd1 _7124_/C sky130_fd_sc_hd__a21o_1
X_8080_ _8080_/A _8080_/B vssd1 vssd1 vccd1 vccd1 _8081_/B sky130_fd_sc_hd__nand2_1
XFILLER_99_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7031_ _6857_/A _7000_/B _7031_/S vssd1 vssd1 vccd1 vccd1 _7032_/B sky130_fd_sc_hd__mux2_1
XFILLER_87_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7933_ _7934_/A _7934_/B vssd1 vssd1 vccd1 vccd1 _8015_/A sky130_fd_sc_hd__or2_1
XFILLER_42_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7864_ _7950_/A _7950_/B vssd1 vssd1 vccd1 vccd1 _7865_/D sky130_fd_sc_hd__nand2_1
XFILLER_51_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6815_ _7007_/B _6853_/A vssd1 vssd1 vccd1 vccd1 _6903_/B sky130_fd_sc_hd__xnor2_1
XFILLER_23_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7795_ _7795_/A _7853_/B vssd1 vssd1 vccd1 vccd1 _7851_/A sky130_fd_sc_hd__xor2_1
X_6746_ _8712_/Q _6746_/B vssd1 vssd1 vccd1 vccd1 _6747_/B sky130_fd_sc_hd__or2_1
XFILLER_51_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6677_ _6677_/A _6677_/B vssd1 vssd1 vccd1 vccd1 _6957_/B sky130_fd_sc_hd__xnor2_2
X_5628_ _5746_/A _5941_/A _6037_/A vssd1 vssd1 vccd1 vccd1 _5628_/X sky130_fd_sc_hd__and3_1
X_8416_ _8461_/B _8414_/A _8461_/A vssd1 vssd1 vccd1 vccd1 _8416_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8347_ _8347_/A _8347_/B vssd1 vssd1 vccd1 vccd1 _8384_/B sky130_fd_sc_hd__xnor2_1
X_5559_ _5559_/A _5559_/B vssd1 vssd1 vccd1 vccd1 _5702_/A sky130_fd_sc_hd__nand2_1
X_8278_ _8278_/A _8250_/B vssd1 vssd1 vccd1 vccd1 _8295_/B sky130_fd_sc_hd__or2b_1
X_7229_ _7232_/A _7232_/B vssd1 vssd1 vccd1 vccd1 _7230_/C sky130_fd_sc_hd__and2_1
XFILLER_86_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_1_0_wb_clk_i clkbuf_3_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_54_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4930_ _4916_/X _4928_/X _4698_/B _5073_/A vssd1 vssd1 vccd1 vccd1 _4930_/X sky130_fd_sc_hd__a211o_1
XFILLER_17_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4861_ _4899_/A _4861_/B _4808_/A vssd1 vssd1 vccd1 vccd1 _4868_/A sky130_fd_sc_hd__or3b_1
XFILLER_45_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6600_ _8712_/Q _6600_/B vssd1 vssd1 vccd1 vccd1 _6747_/A sky130_fd_sc_hd__nand2_1
X_4792_ _6570_/B _4795_/C vssd1 vssd1 vccd1 vccd1 _4822_/B sky130_fd_sc_hd__and2_1
XFILLER_32_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7580_ _7652_/A _7555_/A _7579_/Y _7617_/B vssd1 vssd1 vccd1 vccd1 _7580_/X sky130_fd_sc_hd__a31o_1
X_6531_ _6531_/A _7537_/B _7537_/C vssd1 vssd1 vccd1 vccd1 _6531_/X sky130_fd_sc_hd__and3_1
X_6462_ _8694_/Q _6461_/A _8695_/Q vssd1 vssd1 vccd1 vccd1 _6462_/Y sky130_fd_sc_hd__a21oi_1
X_6393_ _8684_/Q _8688_/Q _8687_/Q _8683_/Q vssd1 vssd1 vccd1 vccd1 _6395_/B sky130_fd_sc_hd__and4bb_1
X_8201_ _8138_/A _8201_/B vssd1 vssd1 vccd1 vccd1 _8201_/X sky130_fd_sc_hd__and2b_1
X_5413_ _5413_/A _5413_/B vssd1 vssd1 vccd1 vccd1 _5415_/A sky130_fd_sc_hd__nor2_1
XFILLER_99_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5344_ _5344_/A _5344_/B vssd1 vssd1 vccd1 vccd1 _8647_/D sky130_fd_sc_hd__nor2_1
X_8132_ _8132_/A _8132_/B vssd1 vssd1 vccd1 vccd1 _8203_/C sky130_fd_sc_hd__xor2_1
XFILLER_87_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5275_ _8727_/Q _5271_/X _5274_/X _5267_/X vssd1 vssd1 vccd1 vccd1 _8628_/D sky130_fd_sc_hd__o211a_1
X_8063_ _8063_/A _8146_/B vssd1 vssd1 vccd1 vccd1 _8309_/A sky130_fd_sc_hd__nand2_1
XFILLER_101_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7014_ _7314_/B _7014_/B vssd1 vssd1 vccd1 vccd1 _7015_/B sky130_fd_sc_hd__and2_1
XFILLER_68_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8896_ _8896_/A _4412_/Y vssd1 vssd1 vccd1 vccd1 io_out[33] sky130_fd_sc_hd__ebufn_8
X_7916_ _8145_/A vssd1 vssd1 vccd1 vccd1 _8308_/A sky130_fd_sc_hd__clkbuf_2
X_7847_ _7847_/A _7847_/B vssd1 vssd1 vccd1 vccd1 _7848_/B sky130_fd_sc_hd__or2_1
XFILLER_62_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7778_ _7885_/A _7972_/A _7777_/X vssd1 vssd1 vccd1 vccd1 _7886_/C sky130_fd_sc_hd__o21a_1
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6729_ _6729_/A _6766_/A vssd1 vssd1 vccd1 vccd1 _7109_/A sky130_fd_sc_hd__xor2_1
XFILLER_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5060_ _5199_/C _5207_/D vssd1 vssd1 vccd1 vccd1 _5231_/B sky130_fd_sc_hd__or2_1
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5962_ _5962_/A _5962_/B vssd1 vssd1 vccd1 vccd1 _6163_/B sky130_fd_sc_hd__xnor2_1
XFILLER_37_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4913_ _5100_/B vssd1 vssd1 vccd1 vccd1 _5107_/C sky130_fd_sc_hd__clkinv_2
X_7701_ _7887_/A vssd1 vssd1 vccd1 vccd1 _7886_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_8681_ _8681_/CLK _8681_/D vssd1 vssd1 vccd1 vccd1 _8681_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5893_ _6118_/A _5893_/B vssd1 vssd1 vccd1 vccd1 _5901_/A sky130_fd_sc_hd__nor2_1
X_4844_ _4844_/A _4919_/A vssd1 vssd1 vccd1 vccd1 _5138_/A sky130_fd_sc_hd__nor2_1
X_7632_ _7908_/A vssd1 vssd1 vccd1 vccd1 _8515_/A sky130_fd_sc_hd__clkbuf_2
X_4775_ _5296_/A vssd1 vssd1 vccd1 vccd1 _7537_/B sky130_fd_sc_hd__buf_2
X_7563_ _8731_/Q _8540_/A _8729_/Q _7562_/Y vssd1 vssd1 vccd1 vccd1 _7563_/X sky130_fd_sc_hd__a31o_1
X_6514_ _6515_/A _6515_/B vssd1 vssd1 vccd1 vccd1 _6516_/A sky130_fd_sc_hd__nor2_1
X_7494_ _7494_/A _7494_/B vssd1 vssd1 vccd1 vccd1 _7501_/B sky130_fd_sc_hd__or2_1
X_6445_ _6446_/B _6446_/C _6444_/Y vssd1 vssd1 vccd1 vccd1 _8688_/D sky130_fd_sc_hd__a21oi_1
X_6376_ _6376_/A _6376_/B vssd1 vssd1 vccd1 vccd1 _8674_/D sky130_fd_sc_hd__nor2_1
X_5327_ _6466_/D _5328_/C _5326_/Y vssd1 vssd1 vccd1 vccd1 _8642_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8115_ _8042_/A _8042_/B _8114_/Y vssd1 vssd1 vccd1 vccd1 _8138_/A sky130_fd_sc_hd__o21a_1
X_8046_ _8046_/A _7975_/B vssd1 vssd1 vccd1 vccd1 _8046_/X sky130_fd_sc_hd__or2b_1
XFILLER_102_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5258_ _5271_/A vssd1 vssd1 vccd1 vccd1 _5258_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_102_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5189_ _5212_/A _5139_/C _5181_/X _5188_/X vssd1 vssd1 vccd1 vccd1 _5190_/C sky130_fd_sc_hd__o31a_1
XFILLER_68_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8879_ _8879_/A _4391_/Y vssd1 vssd1 vccd1 vccd1 io_out[16] sky130_fd_sc_hd__ebufn_8
XFILLER_24_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4560_ _4560_/A vssd1 vssd1 vccd1 vccd1 _8887_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_8_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4491_ _6570_/B vssd1 vssd1 vccd1 vccd1 _4795_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6230_ _6230_/A _6230_/B vssd1 vssd1 vccd1 vccd1 _6283_/B sky130_fd_sc_hd__xor2_4
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6161_ _6012_/B _6161_/B vssd1 vssd1 vccd1 vccd1 _6161_/X sky130_fd_sc_hd__and2b_1
X_5112_ _5243_/A _5136_/B _5067_/Y vssd1 vssd1 vccd1 vccd1 _5112_/X sky130_fd_sc_hd__or3b_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6092_ _6090_/X _6092_/B _6157_/A vssd1 vssd1 vccd1 vccd1 _6094_/A sky130_fd_sc_hd__and3b_1
X_5043_ _5043_/A vssd1 vssd1 vccd1 vccd1 _5143_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_8824__91 vssd1 vssd1 vccd1 vccd1 _8824__91/HI _8933_/A sky130_fd_sc_hd__conb_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6994_ _6991_/Y _6992_/X _6951_/X _6952_/Y vssd1 vssd1 vccd1 vccd1 _7018_/B sky130_fd_sc_hd__o211a_1
XFILLER_92_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8733_ _8733_/CLK _8733_/D vssd1 vssd1 vccd1 vccd1 _8733_/Q sky130_fd_sc_hd__dfxtp_1
X_5945_ _5945_/A _6172_/A vssd1 vssd1 vccd1 vccd1 _5956_/B sky130_fd_sc_hd__xor2_2
XFILLER_80_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5876_ _5713_/X _6070_/B _5876_/S vssd1 vssd1 vccd1 vccd1 _6265_/A sky130_fd_sc_hd__mux2_1
X_8664_ _8732_/CLK _8664_/D vssd1 vssd1 vccd1 vccd1 _8664_/Q sky130_fd_sc_hd__dfxtp_1
X_4827_ _4827_/A _4904_/B vssd1 vssd1 vccd1 vccd1 _5223_/B sky130_fd_sc_hd__nor2_2
X_7615_ _8722_/Q _6423_/X _7614_/X vssd1 vssd1 vccd1 vccd1 _8722_/D sky130_fd_sc_hd__a21bo_1
X_8595_ _8600_/CLK _8595_/D vssd1 vssd1 vccd1 vccd1 _8595_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7546_ _7546_/A _7546_/B vssd1 vssd1 vccd1 vccd1 _7546_/X sky130_fd_sc_hd__or2_1
X_4758_ _4758_/A _4758_/B vssd1 vssd1 vccd1 vccd1 _4844_/A sky130_fd_sc_hd__nand2_2
XFILLER_5_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4689_ _4727_/A _4689_/B _4711_/A vssd1 vssd1 vccd1 vccd1 _4690_/A sky130_fd_sc_hd__and3_1
X_7477_ _7481_/A _7481_/B vssd1 vssd1 vccd1 vccd1 _7482_/A sky130_fd_sc_hd__or2_1
X_6428_ _6432_/C _6428_/B vssd1 vssd1 vccd1 vccd1 _8682_/D sky130_fd_sc_hd__nor2_1
XFILLER_68_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6359_ _6368_/B _6360_/A vssd1 vssd1 vccd1 vccd1 _6366_/A sky130_fd_sc_hd__or2b_1
XFILLER_102_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8029_ _7861_/A _8027_/Y _8028_/X vssd1 vssd1 vccd1 vccd1 _8030_/B sky130_fd_sc_hd__a21o_1
XFILLER_84_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5730_ _5859_/A vssd1 vssd1 vccd1 vccd1 _6030_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_22_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7400_ _7391_/A _7391_/B _7399_/X vssd1 vssd1 vccd1 vccd1 _7467_/A sky130_fd_sc_hd__o21ai_1
XFILLER_30_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5661_ _5661_/A _5661_/B _5661_/C vssd1 vssd1 vccd1 vccd1 _5663_/A sky130_fd_sc_hd__and3_1
X_4612_ _4614_/B _4612_/B _4612_/C vssd1 vssd1 vccd1 vccd1 _4613_/A sky130_fd_sc_hd__and3b_1
X_8380_ _8243_/B _8297_/B _8296_/A vssd1 vssd1 vccd1 vccd1 _8381_/A sky130_fd_sc_hd__a21oi_1
X_5592_ _5661_/A vssd1 vssd1 vccd1 vccd1 _5594_/A sky130_fd_sc_hd__inv_2
X_7331_ _7439_/A _7439_/B vssd1 vssd1 vccd1 vccd1 _7339_/A sky130_fd_sc_hd__xnor2_1
X_4543_ _4567_/B vssd1 vssd1 vccd1 vccd1 _4552_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_7262_ _7260_/A _7260_/B _7267_/B _7267_/A vssd1 vssd1 vccd1 vccd1 _7264_/B sky130_fd_sc_hd__o22a_1
X_4474_ _4720_/A _4714_/A vssd1 vssd1 vccd1 vccd1 _4662_/A sky130_fd_sc_hd__or2_1
X_6213_ _6213_/A _6213_/B vssd1 vssd1 vccd1 vccd1 _6226_/A sky130_fd_sc_hd__xnor2_1
X_7193_ _7193_/A _7193_/B vssd1 vssd1 vccd1 vccd1 _7225_/B sky130_fd_sc_hd__or2_1
X_6144_ _6151_/A _6154_/C vssd1 vssd1 vccd1 vccd1 _6299_/C sky130_fd_sc_hd__or2b_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6075_ _6075_/A _6075_/B vssd1 vssd1 vccd1 vccd1 _6076_/B sky130_fd_sc_hd__nand2_1
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5026_ _5218_/B _5166_/B vssd1 vssd1 vccd1 vccd1 _5027_/C sky130_fd_sc_hd__nor2_1
XFILLER_85_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6977_ _6892_/A _6892_/B _6722_/A _7169_/B vssd1 vssd1 vccd1 vccd1 _6978_/C sky130_fd_sc_hd__a2bb2o_1
XFILLER_26_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8716_ _8734_/CLK _8716_/D vssd1 vssd1 vccd1 vccd1 _8716_/Q sky130_fd_sc_hd__dfxtp_1
X_5928_ _5928_/A _5928_/B vssd1 vssd1 vccd1 vccd1 _6060_/C sky130_fd_sc_hd__xor2_1
X_8647_ _8681_/CLK _8647_/D vssd1 vssd1 vccd1 vccd1 _8647_/Q sky130_fd_sc_hd__dfxtp_1
X_5859_ _5859_/A _5859_/B vssd1 vssd1 vccd1 vccd1 _5941_/C sky130_fd_sc_hd__or2_1
X_8578_ _8578_/A _8578_/B vssd1 vssd1 vccd1 vccd1 _8578_/Y sky130_fd_sc_hd__nor2_1
X_7529_ _7529_/A _7534_/B vssd1 vssd1 vccd1 vccd1 _7529_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_5_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6900_ _6901_/A _6901_/B _6901_/C vssd1 vssd1 vccd1 vccd1 _6902_/A sky130_fd_sc_hd__a21o_1
X_7880_ _7880_/A _7880_/B vssd1 vssd1 vccd1 vccd1 _7881_/C sky130_fd_sc_hd__xor2_1
XFILLER_35_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6831_ _6841_/A _6914_/B vssd1 vssd1 vccd1 vccd1 _6831_/Y sky130_fd_sc_hd__nor2_1
XFILLER_35_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6762_ _6792_/A _6792_/B vssd1 vssd1 vccd1 vccd1 _6763_/B sky130_fd_sc_hd__xnor2_1
XFILLER_23_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8501_ _8501_/A _8501_/B _8510_/A vssd1 vssd1 vccd1 vccd1 _8501_/X sky130_fd_sc_hd__or3_1
X_6693_ _6775_/A vssd1 vssd1 vccd1 vccd1 _6724_/A sky130_fd_sc_hd__clkbuf_2
X_5713_ _5713_/A vssd1 vssd1 vccd1 vccd1 _5713_/X sky130_fd_sc_hd__clkbuf_2
X_5644_ _6028_/A _5952_/B vssd1 vssd1 vccd1 vccd1 _5910_/B sky130_fd_sc_hd__nor2_2
X_8432_ _8433_/A _8433_/B vssd1 vssd1 vccd1 vccd1 _8497_/A sky130_fd_sc_hd__nand2_1
X_8363_ _8166_/X _8289_/A _8288_/B _8362_/X vssd1 vssd1 vccd1 vccd1 _8374_/A sky130_fd_sc_hd__a31o_1
X_7314_ _7314_/A _7314_/B _7314_/C vssd1 vssd1 vccd1 vccd1 _7315_/B sky130_fd_sc_hd__nand3_1
X_5575_ _5575_/A _5788_/B vssd1 vssd1 vccd1 vccd1 _5723_/A sky130_fd_sc_hd__nand2_1
Xclkbuf_4_3_0_wb_clk_i clkbuf_4_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _8671_/CLK
+ sky130_fd_sc_hd__clkbuf_2
X_4526_ _8609_/Q vssd1 vssd1 vccd1 vccd1 _4801_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_8294_ _8295_/A _8295_/B _8295_/C vssd1 vssd1 vccd1 vccd1 _8296_/A sky130_fd_sc_hd__a21oi_1
XFILLER_104_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4457_ _4461_/A vssd1 vssd1 vccd1 vccd1 _4457_/Y sky130_fd_sc_hd__inv_2
X_7245_ _7245_/A _7245_/B _7245_/C vssd1 vssd1 vccd1 vccd1 _7249_/A sky130_fd_sc_hd__nand3_1
XFILLER_49_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7176_ _7182_/A _7182_/B _7175_/Y vssd1 vssd1 vccd1 vccd1 _7178_/A sky130_fd_sc_hd__o21a_1
X_4388_ _4388_/A vssd1 vssd1 vccd1 vccd1 _4388_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6127_ _5560_/A _6071_/C _6136_/A vssd1 vssd1 vccd1 vccd1 _6129_/B sky130_fd_sc_hd__o21a_1
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6058_ _6058_/A _6058_/B vssd1 vssd1 vccd1 vccd1 _6091_/C sky130_fd_sc_hd__xor2_1
X_5009_ _5238_/B _5009_/B _5154_/C _5224_/B vssd1 vssd1 vccd1 vccd1 _5009_/X sky130_fd_sc_hd__or4_1
XFILLER_38_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5360_ _5360_/A vssd1 vssd1 vccd1 vccd1 _8652_/D sky130_fd_sc_hd__clkbuf_1
X_5291_ _8641_/Q _8640_/Q _5289_/X _6466_/D _8643_/Q vssd1 vssd1 vccd1 vccd1 _5291_/X
+ sky130_fd_sc_hd__a311o_1
X_7030_ _7443_/A _6929_/Y _6932_/B _7335_/B vssd1 vssd1 vccd1 vccd1 _7034_/A sky130_fd_sc_hd__a22o_1
XFILLER_101_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7932_ _7818_/A _7817_/B _7817_/A vssd1 vssd1 vccd1 vccd1 _7934_/B sky130_fd_sc_hd__o21ba_1
XFILLER_35_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7863_ _8208_/A _7950_/A _7878_/A vssd1 vssd1 vccd1 vccd1 _7865_/C sky130_fd_sc_hd__a21o_1
X_6814_ _7332_/B _6927_/A vssd1 vssd1 vccd1 vccd1 _6853_/A sky130_fd_sc_hd__nor2_2
XFILLER_50_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7794_ _8515_/D _8122_/B _7794_/C vssd1 vssd1 vccd1 vccd1 _7853_/B sky130_fd_sc_hd__and3_1
X_6745_ _6745_/A _6745_/B vssd1 vssd1 vccd1 vccd1 _6748_/A sky130_fd_sc_hd__nand2_2
X_6676_ _6876_/B _7352_/C vssd1 vssd1 vccd1 vccd1 _6700_/A sky130_fd_sc_hd__nor2_1
X_8415_ _8415_/A _8415_/B _8415_/C vssd1 vssd1 vccd1 vccd1 _8461_/A sky130_fd_sc_hd__and3_1
X_5627_ _5627_/A vssd1 vssd1 vccd1 vccd1 _5941_/A sky130_fd_sc_hd__clkbuf_2
X_8346_ _8346_/A _8346_/B vssd1 vssd1 vccd1 vccd1 _8347_/B sky130_fd_sc_hd__nor2_1
X_5558_ _5533_/A _5558_/B vssd1 vssd1 vccd1 vccd1 _5699_/A sky130_fd_sc_hd__nand2b_1
X_4509_ _4795_/B _4795_/C vssd1 vssd1 vccd1 vccd1 _4820_/B sky130_fd_sc_hd__or2_1
X_8277_ _8277_/A _8277_/B vssd1 vssd1 vccd1 vccd1 _8295_/A sky130_fd_sc_hd__nand2_1
X_7228_ _7228_/A _7228_/B vssd1 vssd1 vccd1 vccd1 _7232_/B sky130_fd_sc_hd__xor2_1
X_5489_ _5374_/A _7871_/A vssd1 vssd1 vccd1 vccd1 _5489_/X sky130_fd_sc_hd__and2b_1
X_7159_ _7159_/A _7159_/B vssd1 vssd1 vccd1 vccd1 _7195_/B sky130_fd_sc_hd__xor2_1
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8785__52 vssd1 vssd1 vccd1 vccd1 _8785__52/HI _8894_/A sky130_fd_sc_hd__conb_1
XFILLER_73_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4860_ _4864_/A _4864_/B vssd1 vssd1 vccd1 vccd1 _4876_/A sky130_fd_sc_hd__nand2_1
XFILLER_17_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6530_ _7548_/B vssd1 vssd1 vccd1 vccd1 _7537_/C sky130_fd_sc_hd__clkbuf_2
X_4791_ _4795_/B _4795_/C vssd1 vssd1 vccd1 vccd1 _4822_/A sky130_fd_sc_hd__nor2_1
XFILLER_20_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6461_ _6461_/A _6461_/B vssd1 vssd1 vccd1 vccd1 _8693_/D sky130_fd_sc_hd__nor2_1
X_6392_ _8678_/Q _8682_/Q _6426_/A _8677_/Q vssd1 vssd1 vccd1 vccd1 _6397_/B sky130_fd_sc_hd__and4bb_1
X_8200_ _8200_/A _8200_/B vssd1 vssd1 vccd1 vccd1 _8240_/A sky130_fd_sc_hd__xor2_1
X_5412_ _8660_/Q _5426_/B vssd1 vssd1 vccd1 vccd1 _5413_/B sky130_fd_sc_hd__and2b_1
X_5343_ _8647_/Q _5345_/C _5323_/X vssd1 vssd1 vccd1 vccd1 _5344_/B sky130_fd_sc_hd__o21ai_1
X_8131_ _8221_/A _8131_/B vssd1 vssd1 vccd1 vccd1 _8132_/B sky130_fd_sc_hd__xnor2_1
XFILLER_99_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5274_ _8628_/Q _5276_/B vssd1 vssd1 vccd1 vccd1 _5274_/X sky130_fd_sc_hd__or2_1
X_8062_ _7905_/B _8065_/B vssd1 vssd1 vccd1 vccd1 _8284_/A sky130_fd_sc_hd__nand2b_2
X_7013_ _7013_/A _7013_/B vssd1 vssd1 vccd1 vccd1 _7014_/B sky130_fd_sc_hd__nand2_1
XFILLER_68_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8895_ _8895_/A _4411_/Y vssd1 vssd1 vccd1 vccd1 io_out[32] sky130_fd_sc_hd__ebufn_8
X_7915_ _8000_/A _8000_/B vssd1 vssd1 vccd1 vccd1 _7922_/A sky130_fd_sc_hd__xnor2_1
XFILLER_36_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7846_ _8102_/A _7846_/B vssd1 vssd1 vccd1 vccd1 _7846_/Y sky130_fd_sc_hd__nand2_1
XFILLER_51_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4989_ _5017_/C vssd1 vssd1 vccd1 vccd1 _5096_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_7777_ _7728_/A _8118_/B _8118_/C _7859_/B _8118_/A vssd1 vssd1 vccd1 vccd1 _7777_/X
+ sky130_fd_sc_hd__a32o_1
X_6728_ _6769_/A _6728_/B vssd1 vssd1 vccd1 vccd1 _6766_/A sky130_fd_sc_hd__xor2_1
XFILLER_11_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6659_ _6659_/A _6659_/B vssd1 vssd1 vccd1 vccd1 _6678_/A sky130_fd_sc_hd__nand2_1
X_8329_ _8228_/A _8338_/B _7963_/X vssd1 vssd1 vccd1 vccd1 _8396_/A sky130_fd_sc_hd__a21o_1
XFILLER_11_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5961_ _5961_/A _5961_/B vssd1 vssd1 vccd1 vccd1 _5962_/B sky130_fd_sc_hd__nor2_1
XFILLER_25_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8680_ _8689_/CLK _8680_/D vssd1 vssd1 vccd1 vccd1 _8680_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4912_ _5047_/A _4876_/A _4872_/X vssd1 vssd1 vccd1 vccd1 _5100_/B sky130_fd_sc_hd__o21a_1
XFILLER_18_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7700_ _7758_/A vssd1 vssd1 vccd1 vccd1 _7887_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7631_ _7722_/A _7722_/B vssd1 vssd1 vccd1 vccd1 _7908_/A sky130_fd_sc_hd__and2_1
X_5892_ _5892_/A vssd1 vssd1 vccd1 vccd1 _6118_/A sky130_fd_sc_hd__clkbuf_2
X_4843_ _4966_/A _5097_/A vssd1 vssd1 vccd1 vccd1 _5127_/A sky130_fd_sc_hd__or2_2
XFILLER_60_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4774_ _4799_/A _4774_/B _4774_/C vssd1 vssd1 vccd1 vccd1 _4781_/B sky130_fd_sc_hd__and3_1
X_7562_ _8563_/A vssd1 vssd1 vccd1 vccd1 _7562_/Y sky130_fd_sc_hd__inv_2
X_6513_ _6509_/A _5362_/X _6508_/X _6512_/X vssd1 vssd1 vccd1 vccd1 _8699_/D sky130_fd_sc_hd__a22o_1
X_7493_ _7493_/A _7493_/B vssd1 vssd1 vccd1 vccd1 _7494_/B sky130_fd_sc_hd__and2_1
XFILLER_20_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6444_ _6446_/B _6446_/C _6406_/B vssd1 vssd1 vccd1 vccd1 _6444_/Y sky130_fd_sc_hd__o21ai_1
X_6375_ _5374_/A _5410_/X _6373_/X _4785_/A vssd1 vssd1 vccd1 vccd1 _6376_/B sky130_fd_sc_hd__a31o_1
X_5326_ _6466_/D _5328_/C _5311_/X vssd1 vssd1 vccd1 vccd1 _5326_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8114_ _8114_/A _8114_/B vssd1 vssd1 vccd1 vccd1 _8114_/Y sky130_fd_sc_hd__nand2_1
X_5257_ _4567_/B _4805_/X _5033_/X _5256_/Y _4765_/B vssd1 vssd1 vccd1 vccd1 _5271_/A
+ sky130_fd_sc_hd__a41o_2
X_8045_ _8045_/A _8045_/B vssd1 vssd1 vccd1 vccd1 _8045_/Y sky130_fd_sc_hd__nand2_1
X_5188_ _5215_/A _5188_/B _5188_/C _5188_/D vssd1 vssd1 vccd1 vccd1 _5188_/X sky130_fd_sc_hd__or4_1
XFILLER_28_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8755__22 vssd1 vssd1 vccd1 vccd1 _8755__22/HI _8850_/A sky130_fd_sc_hd__conb_1
X_8878_ _8878_/A _4390_/Y vssd1 vssd1 vccd1 vccd1 io_out[15] sky130_fd_sc_hd__ebufn_8
XFILLER_24_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7829_ _7850_/A _7850_/B vssd1 vssd1 vccd1 vccd1 _7831_/A sky130_fd_sc_hd__xor2_1
XFILLER_7_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4490_ _8616_/Q vssd1 vssd1 vccd1 vccd1 _6570_/B sky130_fd_sc_hd__buf_4
XFILLER_10_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6160_ _6160_/A _6014_/B vssd1 vssd1 vccd1 vccd1 _6236_/A sky130_fd_sc_hd__or2b_1
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5111_ _5111_/A _5111_/B _5116_/A vssd1 vssd1 vccd1 vccd1 _5136_/C sky130_fd_sc_hd__or3_1
XFILLER_69_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6091_ _6091_/A _6091_/B _6091_/C vssd1 vssd1 vccd1 vccd1 _6092_/B sky130_fd_sc_hd__or3_1
X_5042_ _5143_/A _5208_/A _5078_/C vssd1 vssd1 vccd1 vccd1 _5042_/X sky130_fd_sc_hd__or3_1
XFILLER_84_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6993_ _6951_/X _6952_/Y _6991_/Y _6992_/X vssd1 vssd1 vccd1 vccd1 _7018_/A sky130_fd_sc_hd__a211oi_2
X_5944_ _5944_/A _5944_/B vssd1 vssd1 vccd1 vccd1 _6172_/A sky130_fd_sc_hd__nand2_4
X_8732_ _8732_/CLK _8732_/D vssd1 vssd1 vccd1 vccd1 _8732_/Q sky130_fd_sc_hd__dfxtp_1
X_8663_ _8671_/CLK _8663_/D vssd1 vssd1 vccd1 vccd1 _8663_/Q sky130_fd_sc_hd__dfxtp_1
X_5875_ _5997_/A _6134_/B vssd1 vssd1 vccd1 vccd1 _5876_/S sky130_fd_sc_hd__nor2_1
X_4826_ _4849_/B vssd1 vssd1 vccd1 vccd1 _4904_/B sky130_fd_sc_hd__clkbuf_2
X_8594_ _8600_/CLK _8594_/D vssd1 vssd1 vccd1 vccd1 _8594_/Q sky130_fd_sc_hd__dfxtp_1
X_7614_ _7614_/A _8543_/S _7614_/C _7624_/S vssd1 vssd1 vccd1 vccd1 _7614_/X sky130_fd_sc_hd__or4_1
X_7545_ _7540_/A _7537_/C _7543_/Y _7544_/X vssd1 vssd1 vccd1 vccd1 _8714_/D sky130_fd_sc_hd__a211o_1
X_4757_ _5265_/A vssd1 vssd1 vccd1 vccd1 _5285_/B sky130_fd_sc_hd__clkbuf_2
X_4688_ _4719_/A vssd1 vssd1 vccd1 vccd1 _4711_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7476_ _7479_/B _7475_/C _7475_/A vssd1 vssd1 vccd1 vccd1 _7476_/Y sky130_fd_sc_hd__a21oi_1
X_6427_ _8682_/Q _6425_/A _6406_/B vssd1 vssd1 vccd1 vccd1 _6428_/B sky130_fd_sc_hd__o21ai_1
XFILLER_88_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6358_ _8671_/Q _5410_/X _6356_/Y _6357_/X _4746_/X vssd1 vssd1 vccd1 vccd1 _8671_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_102_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5309_ _8637_/Q _5307_/B _5308_/X vssd1 vssd1 vccd1 vccd1 _5310_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6289_ _6289_/A _6289_/B vssd1 vssd1 vccd1 vccd1 _6290_/B sky130_fd_sc_hd__xnor2_2
X_8028_ _8130_/A _7955_/C _7955_/D _8130_/B _7773_/A vssd1 vssd1 vccd1 vccd1 _8028_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_56_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5660_ _5660_/A _5660_/B vssd1 vssd1 vccd1 vccd1 _5661_/C sky130_fd_sc_hd__nand2_1
XFILLER_90_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4611_ _8588_/Q _4610_/C _8589_/Q vssd1 vssd1 vccd1 vccd1 _4612_/C sky130_fd_sc_hd__a21o_1
X_5591_ _5591_/A _8659_/Q vssd1 vssd1 vccd1 vccd1 _5661_/A sky130_fd_sc_hd__or2b_2
X_7330_ _7003_/A _7003_/B _7329_/X vssd1 vssd1 vccd1 vccd1 _7439_/B sky130_fd_sc_hd__a21oi_2
X_4542_ _4478_/X _4527_/X _4541_/X vssd1 vssd1 vccd1 vccd1 _4567_/B sky130_fd_sc_hd__o21a_2
X_4473_ _6557_/B vssd1 vssd1 vccd1 vccd1 _4714_/A sky130_fd_sc_hd__clkbuf_1
X_7261_ _7280_/B _7261_/B vssd1 vssd1 vccd1 vccd1 _7267_/A sky130_fd_sc_hd__nand2_1
XFILLER_89_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6212_ _5713_/X _5987_/B _6211_/X vssd1 vssd1 vccd1 vccd1 _6213_/B sky130_fd_sc_hd__a21oi_1
X_7192_ _7190_/X _7189_/Y _7188_/Y _7188_/A vssd1 vssd1 vccd1 vccd1 _7193_/B sky130_fd_sc_hd__a211oi_1
XFILLER_97_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6143_ _6143_/A _6143_/B _6143_/C vssd1 vssd1 vccd1 vccd1 _6154_/C sky130_fd_sc_hd__nand3_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6074_ _6075_/A _6075_/B vssd1 vssd1 vccd1 vccd1 _6082_/A sky130_fd_sc_hd__or2_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5025_ _5200_/B vssd1 vssd1 vccd1 vccd1 _5106_/B sky130_fd_sc_hd__clkbuf_2
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6976_ _7366_/B _6975_/C _6975_/A vssd1 vssd1 vccd1 vccd1 _6978_/B sky130_fd_sc_hd__a21o_1
XFILLER_26_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8715_ _8715_/CLK _8715_/D vssd1 vssd1 vccd1 vccd1 _8715_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5927_ _5930_/A _5930_/B vssd1 vssd1 vccd1 vccd1 _5928_/B sky130_fd_sc_hd__xor2_1
XFILLER_41_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8646_ _8677_/CLK _8646_/D vssd1 vssd1 vccd1 vccd1 _8646_/Q sky130_fd_sc_hd__dfxtp_1
X_5858_ _5941_/A vssd1 vssd1 vccd1 vccd1 _6119_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4809_ _4879_/A vssd1 vssd1 vccd1 vccd1 _4885_/B sky130_fd_sc_hd__clkbuf_2
X_8577_ _8572_/A _8576_/X _8577_/S vssd1 vssd1 vccd1 vccd1 _8578_/B sky130_fd_sc_hd__mux2_1
X_5789_ _5798_/A _6211_/B _6221_/A vssd1 vssd1 vccd1 vccd1 _5790_/B sky130_fd_sc_hd__o21ai_1
X_7528_ _7523_/A _7523_/B _7521_/A vssd1 vssd1 vccd1 vccd1 _7534_/B sky130_fd_sc_hd__a21oi_1
XFILLER_5_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7459_ _7459_/A _7459_/B vssd1 vssd1 vccd1 vccd1 _7460_/B sky130_fd_sc_hd__xor2_1
XFILLER_79_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6830_ _6931_/B vssd1 vssd1 vccd1 vccd1 _6914_/B sky130_fd_sc_hd__buf_2
XFILLER_90_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6761_ _6793_/C _7127_/A _7103_/A vssd1 vssd1 vccd1 vccd1 _6792_/B sky130_fd_sc_hd__a21oi_1
XFILLER_62_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5712_ _5775_/A _5775_/B vssd1 vssd1 vccd1 vccd1 _5720_/A sky130_fd_sc_hd__xnor2_1
X_8500_ _8509_/B _8509_/C _8509_/A vssd1 vssd1 vccd1 vccd1 _8510_/A sky130_fd_sc_hd__a21oi_1
X_6692_ _7254_/A _6890_/A vssd1 vssd1 vccd1 vccd1 _6775_/A sky130_fd_sc_hd__nor2_1
XFILLER_31_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8431_ _8431_/A _8431_/B vssd1 vssd1 vccd1 vccd1 _8433_/B sky130_fd_sc_hd__xnor2_1
X_5643_ _5609_/B _5614_/B _5634_/X vssd1 vssd1 vccd1 vccd1 _5952_/B sky130_fd_sc_hd__a21o_1
X_8362_ _8290_/A _8362_/B vssd1 vssd1 vccd1 vccd1 _8362_/X sky130_fd_sc_hd__and2b_1
X_5574_ _5574_/A vssd1 vssd1 vccd1 vccd1 _5788_/B sky130_fd_sc_hd__buf_2
X_7313_ _7314_/A _7314_/B _7314_/C vssd1 vssd1 vccd1 vccd1 _7315_/A sky130_fd_sc_hd__a21o_1
X_4525_ _6605_/B vssd1 vssd1 vccd1 vccd1 _4733_/S sky130_fd_sc_hd__dlymetal6s2s_1
X_8293_ _8375_/B _8293_/B vssd1 vssd1 vccd1 vccd1 _8295_/C sky130_fd_sc_hd__xor2_1
X_4456_ _4456_/A vssd1 vssd1 vccd1 vccd1 _4461_/A sky130_fd_sc_hd__clkbuf_4
X_7244_ _7223_/A _7223_/C _7223_/B vssd1 vssd1 vccd1 vccd1 _7245_/C sky130_fd_sc_hd__o21ai_1
X_4387_ _4388_/A vssd1 vssd1 vccd1 vccd1 _4387_/Y sky130_fd_sc_hd__inv_2
X_7175_ _7234_/A _7175_/B vssd1 vssd1 vccd1 vccd1 _7175_/Y sky130_fd_sc_hd__nand2_1
XFILLER_58_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6126_ _6126_/A _6126_/B _6126_/C vssd1 vssd1 vccd1 vccd1 _6136_/A sky130_fd_sc_hd__or3_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6057_ _6089_/A _6089_/B vssd1 vssd1 vccd1 vccd1 _6091_/B sky130_fd_sc_hd__and2_1
XFILLER_45_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5008_ _5233_/B _5054_/A vssd1 vssd1 vccd1 vccd1 _5224_/B sky130_fd_sc_hd__or2_2
X_6959_ _6958_/B _6958_/C _6892_/B vssd1 vssd1 vccd1 vccd1 _6960_/C sky130_fd_sc_hd__o21ai_1
X_8629_ _8734_/CLK _8629_/D vssd1 vssd1 vccd1 vccd1 _8629_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5290_ _8642_/Q vssd1 vssd1 vccd1 vccd1 _6466_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_4_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7931_ _7928_/X _7929_/Y _7851_/X _7852_/Y vssd1 vssd1 vccd1 vccd1 _7936_/B sky130_fd_sc_hd__o211a_1
XFILLER_82_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7862_ _7862_/A _8130_/A vssd1 vssd1 vccd1 vccd1 _7878_/A sky130_fd_sc_hd__nor2_1
X_6813_ _6813_/A vssd1 vssd1 vccd1 vccd1 _6927_/A sky130_fd_sc_hd__buf_2
XFILLER_50_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7793_ _7885_/A _8124_/A vssd1 vssd1 vccd1 vccd1 _7794_/C sky130_fd_sc_hd__nand2_1
X_6744_ _6744_/A vssd1 vssd1 vccd1 vccd1 _7010_/A sky130_fd_sc_hd__clkbuf_2
X_6675_ _7074_/C vssd1 vssd1 vccd1 vccd1 _7352_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_5626_ _5742_/A vssd1 vssd1 vccd1 vccd1 _5746_/A sky130_fd_sc_hd__clkbuf_2
X_8414_ _8414_/A _8414_/B vssd1 vssd1 vccd1 vccd1 _8461_/B sky130_fd_sc_hd__nor2_1
X_8345_ _8345_/A _8345_/B _8345_/C vssd1 vssd1 vccd1 vccd1 _8346_/B sky130_fd_sc_hd__and3_1
X_5557_ _5550_/A _5557_/B vssd1 vssd1 vccd1 vccd1 _5583_/A sky130_fd_sc_hd__and2b_1
XFILLER_104_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4508_ _8614_/Q _8613_/Q _7630_/B vssd1 vssd1 vccd1 vccd1 _4795_/C sky130_fd_sc_hd__o21a_1
X_8276_ _8199_/A _8199_/B _8200_/B _8200_/A vssd1 vssd1 vccd1 vccd1 _8298_/A sky130_fd_sc_hd__o2bb2a_1
X_5488_ _5540_/A _5527_/B vssd1 vssd1 vccd1 vccd1 _5502_/A sky130_fd_sc_hd__nand2_1
X_7227_ _7010_/B _6914_/B _7146_/B _7465_/A vssd1 vssd1 vccd1 vccd1 _7232_/A sky130_fd_sc_hd__o22ai_4
X_4439_ _4443_/A vssd1 vssd1 vccd1 vccd1 _4439_/Y sky130_fd_sc_hd__inv_2
X_7158_ _7152_/A _7152_/B _7157_/X vssd1 vssd1 vccd1 vccd1 _7195_/A sky130_fd_sc_hd__o21a_1
X_7089_ _7135_/A _7135_/B vssd1 vssd1 vccd1 vccd1 _7089_/Y sky130_fd_sc_hd__nand2_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6109_ _6116_/A _6116_/B vssd1 vssd1 vccd1 vccd1 _6117_/A sky130_fd_sc_hd__or2_1
XFILLER_46_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4790_ _4790_/A vssd1 vssd1 vccd1 vccd1 _4790_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6460_ _8693_/Q _6459_/B _6401_/B vssd1 vssd1 vccd1 vccd1 _6461_/B sky130_fd_sc_hd__o21ai_1
XFILLER_9_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6391_ _8676_/Q _8675_/Q vssd1 vssd1 vccd1 vccd1 _6397_/A sky130_fd_sc_hd__nor2_1
X_5411_ _5425_/B _5411_/B vssd1 vssd1 vccd1 vccd1 _5413_/A sky130_fd_sc_hd__and2b_1
X_5342_ _8647_/Q _5345_/C vssd1 vssd1 vccd1 vccd1 _5344_/A sky130_fd_sc_hd__and2_1
X_8130_ _8130_/A _8130_/B vssd1 vssd1 vccd1 vccd1 _8221_/A sky130_fd_sc_hd__or2_2
X_8061_ _8061_/A _8489_/A vssd1 vssd1 vccd1 vccd1 _8076_/C sky130_fd_sc_hd__xnor2_1
X_7012_ _7013_/A _7013_/B vssd1 vssd1 vccd1 vccd1 _7314_/B sky130_fd_sc_hd__or2_1
X_5273_ _8726_/Q _5271_/X _5272_/X _5267_/X vssd1 vssd1 vccd1 vccd1 _8627_/D sky130_fd_sc_hd__o211a_1
XFILLER_99_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8894_ _8894_/A _4410_/Y vssd1 vssd1 vccd1 vccd1 io_out[31] sky130_fd_sc_hd__ebufn_8
X_7914_ _7914_/A _7984_/B vssd1 vssd1 vccd1 vccd1 _8000_/B sky130_fd_sc_hd__xnor2_1
XFILLER_62_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7845_ _8533_/A _7848_/A vssd1 vssd1 vccd1 vccd1 _7846_/B sky130_fd_sc_hd__nand2_1
XFILLER_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4988_ _5190_/A _4970_/B _4985_/X _4987_/X _4711_/B vssd1 vssd1 vccd1 vccd1 _4988_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_23_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7776_ _7771_/A _7771_/C _7771_/B vssd1 vssd1 vccd1 vccd1 _8118_/C sky130_fd_sc_hd__a21o_1
X_6727_ _6727_/A _6795_/A vssd1 vssd1 vccd1 vccd1 _6728_/B sky130_fd_sc_hd__xnor2_1
X_6658_ _6688_/A _6689_/A _6657_/A vssd1 vssd1 vccd1 vccd1 _7074_/C sky130_fd_sc_hd__a21oi_4
X_5609_ _5732_/A _5609_/B vssd1 vssd1 vccd1 vccd1 _5641_/A sky130_fd_sc_hd__nand2_1
X_6589_ _6589_/A vssd1 vssd1 vccd1 vccd1 _7454_/A sky130_fd_sc_hd__buf_2
XFILLER_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8328_ _8328_/A _8328_/B vssd1 vssd1 vccd1 vccd1 _8345_/A sky130_fd_sc_hd__or2_1
XFILLER_87_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8259_ _8259_/A _8259_/B vssd1 vssd1 vccd1 vccd1 _8260_/B sky130_fd_sc_hd__xnor2_2
XFILLER_78_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5960_ _5960_/A _5960_/B _5960_/C vssd1 vssd1 vccd1 vccd1 _5961_/B sky130_fd_sc_hd__and3_1
X_4911_ _5154_/B vssd1 vssd1 vccd1 vccd1 _5017_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_18_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5891_ _5891_/A _5891_/B vssd1 vssd1 vccd1 vccd1 _5903_/A sky130_fd_sc_hd__xnor2_2
XFILLER_33_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7630_ _7630_/A _7630_/B vssd1 vssd1 vccd1 vccd1 _7722_/B sky130_fd_sc_hd__nand2_1
X_4842_ _4998_/B _5222_/D vssd1 vssd1 vccd1 vccd1 _5097_/A sky130_fd_sc_hd__or2_1
XFILLER_21_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4773_ _4774_/B _4779_/B _4772_/Y vssd1 vssd1 vccd1 vccd1 _8617_/D sky130_fd_sc_hd__a21oi_1
X_7561_ _8553_/A _8571_/B vssd1 vssd1 vccd1 vccd1 _8563_/A sky130_fd_sc_hd__and2_1
XFILLER_20_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6512_ _6510_/Y _6512_/B vssd1 vssd1 vccd1 vccd1 _6512_/X sky130_fd_sc_hd__and2b_1
X_7492_ _7501_/A _7510_/A vssd1 vssd1 vccd1 vccd1 _7492_/X sky130_fd_sc_hd__and2b_1
X_6443_ _6446_/C _6443_/B vssd1 vssd1 vccd1 vccd1 _8687_/D sky130_fd_sc_hd__nor2_1
X_6374_ _5410_/X _6373_/X _5374_/A vssd1 vssd1 vccd1 vccd1 _6376_/A sky130_fd_sc_hd__a21oi_1
X_5325_ _5328_/C _5325_/B vssd1 vssd1 vccd1 vccd1 _8641_/D sky130_fd_sc_hd__nor2_1
X_8113_ _8049_/A _8049_/B _8112_/X vssd1 vssd1 vccd1 vccd1 _8192_/A sky130_fd_sc_hd__a21oi_2
XFILLER_102_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5256_ _5256_/A _5256_/B vssd1 vssd1 vccd1 vccd1 _5256_/Y sky130_fd_sc_hd__nand2_1
X_8044_ _8044_/A vssd1 vssd1 vccd1 vccd1 _8139_/B sky130_fd_sc_hd__buf_2
X_5187_ _5186_/A _5227_/B _5183_/X _5186_/X vssd1 vssd1 vccd1 vccd1 _5188_/D sky130_fd_sc_hd__o31a_1
XFILLER_28_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8877_ _8877_/A _4388_/Y vssd1 vssd1 vccd1 vccd1 io_out[14] sky130_fd_sc_hd__ebufn_8
XFILLER_24_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7828_ _7940_/A _7828_/B vssd1 vssd1 vccd1 vccd1 _7850_/B sky130_fd_sc_hd__nand2_1
X_8770__37 vssd1 vssd1 vccd1 vccd1 _8770__37/HI _8865_/A sky130_fd_sc_hd__conb_1
X_7759_ _7759_/A _7759_/B vssd1 vssd1 vccd1 vccd1 _7862_/A sky130_fd_sc_hd__xnor2_1
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5110_ _5155_/A _5106_/X _5109_/X _5017_/C vssd1 vssd1 vccd1 vccd1 _5110_/X sky130_fd_sc_hd__a211o_1
XFILLER_88_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6090_ _6152_/A _6152_/B vssd1 vssd1 vccd1 vccd1 _6090_/X sky130_fd_sc_hd__or2b_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5041_ _5050_/C vssd1 vssd1 vccd1 vccd1 _5078_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
XFILLER_65_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6992_ _7347_/A _7347_/B _7347_/C _7347_/D vssd1 vssd1 vccd1 vccd1 _6992_/X sky130_fd_sc_hd__o22a_1
XFILLER_53_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8731_ _8732_/CLK _8731_/D vssd1 vssd1 vccd1 vccd1 _8731_/Q sky130_fd_sc_hd__dfxtp_1
X_5943_ _5943_/A _5952_/B vssd1 vssd1 vccd1 vccd1 _5973_/A sky130_fd_sc_hd__nor2_2
XFILLER_80_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5874_ _5874_/A _5874_/B vssd1 vssd1 vccd1 vccd1 _6134_/B sky130_fd_sc_hd__xnor2_4
X_8662_ _8674_/CLK _8662_/D vssd1 vssd1 vccd1 vccd1 _8662_/Q sky130_fd_sc_hd__dfxtp_1
X_4825_ _4837_/B vssd1 vssd1 vccd1 vccd1 _4849_/B sky130_fd_sc_hd__clkbuf_2
X_8593_ _8600_/CLK _8593_/D vssd1 vssd1 vccd1 vccd1 _8593_/Q sky130_fd_sc_hd__dfxtp_1
X_7613_ _7613_/A _7613_/B _7613_/C vssd1 vssd1 vccd1 vccd1 _7624_/S sky130_fd_sc_hd__and3_1
X_7544_ _7614_/A vssd1 vssd1 vccd1 vccd1 _7544_/X sky130_fd_sc_hd__buf_2
XFILLER_21_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4756_ _7499_/A vssd1 vssd1 vccd1 vccd1 _8544_/A sky130_fd_sc_hd__buf_2
X_4687_ _4763_/A _4687_/B vssd1 vssd1 vccd1 vccd1 _4719_/A sky130_fd_sc_hd__nand2_1
X_7475_ _7475_/A _7479_/B _7475_/C vssd1 vssd1 vccd1 vccd1 _7475_/X sky130_fd_sc_hd__and3_1
X_6426_ _6426_/A _8682_/Q _6426_/C vssd1 vssd1 vccd1 vccd1 _6432_/C sky130_fd_sc_hd__and3_1
X_6357_ _6356_/A _6356_/B _4581_/B vssd1 vssd1 vccd1 vccd1 _6357_/X sky130_fd_sc_hd__a21o_1
XFILLER_102_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5308_ _5323_/A vssd1 vssd1 vccd1 vccd1 _5308_/X sky130_fd_sc_hd__buf_2
XFILLER_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6288_ _6288_/A _6288_/B vssd1 vssd1 vccd1 vccd1 _6289_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5239_ _5218_/B _5128_/B _5243_/B _5237_/A vssd1 vssd1 vccd1 vccd1 _5239_/X sky130_fd_sc_hd__o31a_1
X_8815__82 vssd1 vssd1 vccd1 vccd1 _8815__82/HI _8924_/A sky130_fd_sc_hd__conb_1
XFILLER_29_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8027_ _8122_/C _8130_/B vssd1 vssd1 vccd1 vccd1 _8027_/Y sky130_fd_sc_hd__nor2_1
XFILLER_29_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8929_ _8929_/A _4449_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[28] sky130_fd_sc_hd__ebufn_8
XFILLER_12_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4610_ _8588_/Q _8589_/Q _4610_/C vssd1 vssd1 vccd1 vccd1 _4614_/B sky130_fd_sc_hd__and3_1
X_5590_ _5642_/A _5638_/B _5589_/X vssd1 vssd1 vccd1 vccd1 _5595_/A sky130_fd_sc_hd__a21oi_2
X_4541_ _4541_/A _4541_/B _4668_/A _4541_/D vssd1 vssd1 vccd1 vccd1 _4541_/X sky130_fd_sc_hd__and4_1
X_7260_ _7260_/A _7260_/B vssd1 vssd1 vccd1 vccd1 _7267_/B sky130_fd_sc_hd__xnor2_1
X_4472_ _8607_/Q vssd1 vssd1 vccd1 vccd1 _6557_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_104_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7191_ _7188_/A _7188_/Y _7189_/Y _7190_/X vssd1 vssd1 vccd1 vccd1 _7193_/A sky130_fd_sc_hd__o211a_1
X_6211_ _5986_/B _6211_/B vssd1 vssd1 vccd1 vccd1 _6211_/X sky130_fd_sc_hd__and2b_1
X_6142_ _6143_/A _6143_/B _6143_/C vssd1 vssd1 vccd1 vccd1 _6151_/A sky130_fd_sc_hd__a21oi_2
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6073_ _6073_/A _6073_/B vssd1 vssd1 vccd1 vccd1 _6110_/A sky130_fd_sc_hd__xnor2_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5024_ _4694_/A _5096_/B _5010_/X _5023_/X _4697_/X vssd1 vssd1 vccd1 vccd1 _5024_/X
+ sky130_fd_sc_hd__o32a_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6975_ _6975_/A _7366_/B _6975_/C vssd1 vssd1 vccd1 vccd1 _6978_/A sky130_fd_sc_hd__nand3_1
XFILLER_53_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8714_ _8714_/CLK _8714_/D vssd1 vssd1 vccd1 vccd1 _8714_/Q sky130_fd_sc_hd__dfxtp_1
X_5926_ _5926_/A _5926_/B vssd1 vssd1 vccd1 vccd1 _5930_/B sky130_fd_sc_hd__xnor2_1
X_8645_ _8681_/CLK _8645_/D vssd1 vssd1 vccd1 vccd1 _8645_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5857_ _5829_/A _5829_/B _5856_/Y vssd1 vssd1 vccd1 vccd1 _5933_/A sky130_fd_sc_hd__a21oi_1
X_4808_ _4808_/A _4822_/A _4822_/B _4861_/B vssd1 vssd1 vccd1 vccd1 _4879_/A sky130_fd_sc_hd__or4b_4
X_8576_ _8576_/A _8576_/B vssd1 vssd1 vccd1 vccd1 _8576_/X sky130_fd_sc_hd__or2_1
XFILLER_21_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5788_ _5788_/A _5788_/B vssd1 vssd1 vccd1 vccd1 _6221_/A sky130_fd_sc_hd__nand2_2
X_7527_ _7535_/A _7527_/B vssd1 vssd1 vccd1 vccd1 _7529_/A sky130_fd_sc_hd__nor2_1
X_4739_ _4891_/A _4752_/A vssd1 vssd1 vccd1 vccd1 _4740_/B sky130_fd_sc_hd__nor2_1
X_7458_ _7458_/A _7458_/B vssd1 vssd1 vccd1 vccd1 _7459_/B sky130_fd_sc_hd__xnor2_1
X_6409_ _8676_/Q _8675_/Q _8677_/Q vssd1 vssd1 vccd1 vccd1 _6410_/B sky130_fd_sc_hd__a21o_1
X_7389_ _7463_/A _7463_/B vssd1 vssd1 vccd1 vccd1 _7390_/B sky130_fd_sc_hd__xnor2_1
XFILLER_88_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6760_ _6803_/B _6804_/C vssd1 vssd1 vccd1 vccd1 _6792_/A sky130_fd_sc_hd__xor2_2
X_5711_ _5987_/A _5711_/B vssd1 vssd1 vccd1 vccd1 _5775_/B sky130_fd_sc_hd__xnor2_1
X_6691_ _6625_/X _6688_/X _6689_/X _6876_/A vssd1 vssd1 vccd1 vccd1 _6890_/A sky130_fd_sc_hd__a31o_1
X_8430_ _8430_/A _8430_/B vssd1 vssd1 vccd1 vccd1 _8433_/A sky130_fd_sc_hd__or2_1
X_5642_ _5642_/A _5642_/B vssd1 vssd1 vccd1 vccd1 _6028_/A sky130_fd_sc_hd__and2_2
X_8361_ _8316_/A _8316_/B _8317_/B _8317_/A vssd1 vssd1 vccd1 vccd1 _8439_/B sky130_fd_sc_hd__a2bb2o_1
X_5573_ _5699_/A _5699_/B vssd1 vssd1 vccd1 vccd1 _5582_/A sky130_fd_sc_hd__xnor2_1
X_7312_ _7312_/A _7312_/B vssd1 vssd1 vccd1 vccd1 _7314_/C sky130_fd_sc_hd__xnor2_1
X_4524_ _5190_/A _4986_/B vssd1 vssd1 vccd1 vccd1 _4524_/X sky130_fd_sc_hd__or2_1
X_8292_ _8292_/A _8292_/B vssd1 vssd1 vccd1 vccd1 _8293_/B sky130_fd_sc_hd__xnor2_1
XFILLER_104_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4455_ _4455_/A vssd1 vssd1 vccd1 vccd1 _4455_/Y sky130_fd_sc_hd__inv_2
X_7243_ _7252_/B _7252_/A vssd1 vssd1 vccd1 vccd1 _7245_/B sky130_fd_sc_hd__and2b_1
X_4386_ _4388_/A vssd1 vssd1 vccd1 vccd1 _4386_/Y sky130_fd_sc_hd__inv_2
X_7174_ _7234_/A _7175_/B vssd1 vssd1 vccd1 vccd1 _7182_/B sky130_fd_sc_hd__xnor2_1
XFILLER_98_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6125_ _6020_/B _5567_/B _6071_/A _5981_/A vssd1 vssd1 vccd1 vccd1 _6126_/C sky130_fd_sc_hd__o2bb2a_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6056_ _6056_/A _6056_/B vssd1 vssd1 vccd1 vccd1 _6089_/B sky130_fd_sc_hd__xnor2_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5007_ _5007_/A _5007_/B vssd1 vssd1 vccd1 vccd1 _5154_/C sky130_fd_sc_hd__or2_1
XFILLER_54_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6958_ _6958_/A _6958_/B _6958_/C vssd1 vssd1 vccd1 vccd1 _6960_/B sky130_fd_sc_hd__or3_1
XFILLER_53_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6889_ _7003_/A _6889_/B vssd1 vssd1 vccd1 vccd1 _6897_/A sky130_fd_sc_hd__xnor2_1
X_5909_ _6182_/A _5909_/B vssd1 vssd1 vccd1 vccd1 _5937_/A sky130_fd_sc_hd__nand2_1
X_8628_ _8734_/CLK _8628_/D vssd1 vssd1 vccd1 vccd1 _8628_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8559_ _8560_/B _8576_/A vssd1 vssd1 vccd1 vccd1 _8569_/A sky130_fd_sc_hd__and2b_1
XFILLER_5_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7930_ _7851_/X _7852_/Y _7928_/X _7929_/Y vssd1 vssd1 vccd1 vccd1 _7936_/A sky130_fd_sc_hd__a211oi_2
XFILLER_48_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7861_ _7861_/A vssd1 vssd1 vccd1 vccd1 _7887_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6812_ _6812_/A _6812_/B vssd1 vssd1 vccd1 vccd1 _6813_/A sky130_fd_sc_hd__xnor2_2
XFILLER_23_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7792_ _7792_/A _7792_/B vssd1 vssd1 vccd1 vccd1 _7795_/A sky130_fd_sc_hd__xnor2_1
X_6743_ _7091_/A _7091_/B _6742_/Y vssd1 vssd1 vccd1 vccd1 _6765_/A sky130_fd_sc_hd__a21o_1
X_6674_ _7074_/B vssd1 vssd1 vccd1 vccd1 _6876_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_5625_ _5813_/A vssd1 vssd1 vccd1 vccd1 _5742_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_8413_ _8415_/A _8413_/B vssd1 vssd1 vccd1 vccd1 _8414_/B sky130_fd_sc_hd__nor2_1
X_8344_ _8345_/A _8345_/B _8345_/C vssd1 vssd1 vccd1 vccd1 _8346_/A sky130_fd_sc_hd__a21oi_1
X_5556_ _5556_/A _6024_/A vssd1 vssd1 vccd1 vccd1 _5694_/A sky130_fd_sc_hd__nand2_1
X_4507_ _8615_/Q vssd1 vssd1 vccd1 vccd1 _7630_/B sky130_fd_sc_hd__clkbuf_4
X_8275_ _8260_/A _8260_/B _8274_/Y vssd1 vssd1 vccd1 vccd1 _8355_/B sky130_fd_sc_hd__a21o_1
X_5487_ _6338_/S _8605_/Q vssd1 vssd1 vccd1 vccd1 _5527_/B sky130_fd_sc_hd__nand2_1
XFILLER_104_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4438_ _4456_/A vssd1 vssd1 vccd1 vccd1 _4443_/A sky130_fd_sc_hd__clkbuf_2
X_7226_ _7228_/A _7228_/B vssd1 vssd1 vccd1 vccd1 _7230_/B sky130_fd_sc_hd__nor2_1
XFILLER_98_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4369_ _4369_/A vssd1 vssd1 vccd1 vccd1 _4369_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7157_ _7157_/A _7157_/B vssd1 vssd1 vccd1 vccd1 _7157_/X sky130_fd_sc_hd__or2_1
XFILLER_58_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7088_ _7133_/A _7088_/B vssd1 vssd1 vccd1 vccd1 _7136_/B sky130_fd_sc_hd__xor2_2
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6108_ _6108_/A _6108_/B vssd1 vssd1 vccd1 vccd1 _6116_/B sky130_fd_sc_hd__xnor2_1
XFILLER_100_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6039_ _6039_/A _6039_/B vssd1 vssd1 vccd1 vccd1 _6063_/B sky130_fd_sc_hd__xnor2_1
XFILLER_54_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8776__43 vssd1 vssd1 vccd1 vccd1 _8776__43/HI _8871_/A sky130_fd_sc_hd__conb_1
XFILLER_17_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6390_ _8695_/Q _6390_/B vssd1 vssd1 vccd1 vccd1 _6403_/B sky130_fd_sc_hd__nand2_1
X_5410_ _5410_/A vssd1 vssd1 vccd1 vccd1 _5410_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_99_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5341_ _5341_/A vssd1 vssd1 vccd1 vccd1 _8646_/D sky130_fd_sc_hd__clkbuf_1
X_8060_ _8060_/A vssd1 vssd1 vccd1 vccd1 _8489_/A sky130_fd_sc_hd__clkbuf_2
X_7011_ _6619_/Y _7416_/A _7314_/A vssd1 vssd1 vccd1 vccd1 _7013_/B sky130_fd_sc_hd__a21bo_1
X_5272_ _8627_/Q _5276_/B vssd1 vssd1 vccd1 vccd1 _5272_/X sky130_fd_sc_hd__or2_1
XFILLER_95_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7913_ _7919_/A _7985_/B vssd1 vssd1 vccd1 vccd1 _7984_/B sky130_fd_sc_hd__xnor2_1
X_8893_ _8893_/A _4409_/Y vssd1 vssd1 vccd1 vccd1 io_out[30] sky130_fd_sc_hd__ebufn_8
XFILLER_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7844_ _8533_/A _7848_/A vssd1 vssd1 vccd1 vccd1 _8102_/A sky130_fd_sc_hd__or2_1
XFILLER_36_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7775_ _7775_/A _7775_/B _7771_/B vssd1 vssd1 vccd1 vccd1 _8118_/B sky130_fd_sc_hd__or3b_1
X_6726_ _6697_/B _6697_/C _6697_/A vssd1 vssd1 vccd1 vccd1 _6795_/A sky130_fd_sc_hd__a21boi_2
X_4987_ _5166_/B _4987_/B _4987_/C _4987_/D vssd1 vssd1 vccd1 vccd1 _4987_/X sky130_fd_sc_hd__or4_1
XFILLER_51_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6657_ _6657_/A _6688_/A _6689_/A vssd1 vssd1 vccd1 vccd1 _7074_/B sky130_fd_sc_hd__and3_1
X_6588_ _6588_/A _6588_/B vssd1 vssd1 vccd1 vccd1 _6589_/A sky130_fd_sc_hd__nand2_1
X_5608_ _5634_/A _7906_/B vssd1 vssd1 vccd1 vccd1 _5609_/B sky130_fd_sc_hd__or2_1
XFILLER_3_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8327_ _8388_/A _8327_/B vssd1 vssd1 vccd1 vccd1 _8347_/A sky130_fd_sc_hd__xnor2_1
X_5539_ _6020_/A _5792_/B _5539_/C vssd1 vssd1 vccd1 vccd1 _5548_/B sky130_fd_sc_hd__and3_1
X_8258_ _8258_/A _8258_/B vssd1 vssd1 vccd1 vccd1 _8259_/B sky130_fd_sc_hd__nand2_2
X_7209_ _7210_/A _7210_/B vssd1 vssd1 vccd1 vccd1 _7209_/X sky130_fd_sc_hd__or2b_1
X_8189_ _8180_/A _8180_/B _8179_/A vssd1 vssd1 vccd1 vccd1 _8262_/A sky130_fd_sc_hd__o21ai_2
XFILLER_59_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4910_ _5038_/A _4991_/B _5220_/B vssd1 vssd1 vccd1 vccd1 _5154_/B sky130_fd_sc_hd__nor3_2
X_5890_ _5983_/A _5983_/B vssd1 vssd1 vccd1 vccd1 _5891_/B sky130_fd_sc_hd__xnor2_1
XFILLER_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4841_ _5054_/A _4999_/A vssd1 vssd1 vccd1 vccd1 _5222_/D sky130_fd_sc_hd__or2_1
XFILLER_45_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4772_ _4774_/B _4779_/B _4771_/X vssd1 vssd1 vccd1 vccd1 _4772_/Y sky130_fd_sc_hd__o21ai_1
X_7560_ _8560_/B vssd1 vssd1 vccd1 vccd1 _8571_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6511_ _6565_/A _6511_/B vssd1 vssd1 vccd1 vccd1 _6512_/B sky130_fd_sc_hd__nand2_1
X_7491_ _7491_/A _7491_/B _7491_/C _7491_/D vssd1 vssd1 vccd1 vccd1 _7510_/A sky130_fd_sc_hd__and4_1
X_6442_ _8687_/Q _6441_/B _6423_/X vssd1 vssd1 vccd1 vccd1 _6443_/B sky130_fd_sc_hd__o21ai_1
X_8112_ _8043_/B _8112_/B vssd1 vssd1 vccd1 vccd1 _8112_/X sky130_fd_sc_hd__and2b_1
Xclkbuf_3_0_0_wb_clk_i clkbuf_3_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
X_6373_ _6369_/A _6372_/X _6373_/S vssd1 vssd1 vccd1 vccd1 _6373_/X sky130_fd_sc_hd__mux2_1
X_5324_ _8641_/Q _5321_/A _5323_/X vssd1 vssd1 vccd1 vccd1 _5325_/B sky130_fd_sc_hd__o21ai_1
XFILLER_87_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5255_ _5149_/X _5253_/X _5255_/S vssd1 vssd1 vccd1 vccd1 _5256_/B sky130_fd_sc_hd__mux2_1
X_8043_ _8112_/B _8043_/B vssd1 vssd1 vccd1 vccd1 _8049_/A sky130_fd_sc_hd__xnor2_2
X_5186_ _5186_/A _5223_/A _5186_/C _5186_/D vssd1 vssd1 vccd1 vccd1 _5186_/X sky130_fd_sc_hd__or4_1
XFILLER_68_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8876_ _8876_/A _4387_/Y vssd1 vssd1 vccd1 vccd1 io_out[13] sky130_fd_sc_hd__ebufn_8
X_7827_ _7852_/A _7826_/C _7826_/A vssd1 vssd1 vccd1 vccd1 _7828_/B sky130_fd_sc_hd__o21ai_1
XFILLER_11_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7758_ _7758_/A _7785_/A vssd1 vssd1 vccd1 vccd1 _7779_/A sky130_fd_sc_hd__nand2_1
XFILLER_11_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6709_ _6625_/X _6688_/X _6689_/X _6876_/A _7075_/A vssd1 vssd1 vccd1 vccd1 _6774_/S
+ sky130_fd_sc_hd__a311o_4
X_7689_ _7689_/A _7689_/B vssd1 vssd1 vccd1 vccd1 _7713_/B sky130_fd_sc_hd__nor2_4
XFILLER_78_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8746__13 vssd1 vssd1 vccd1 vccd1 _8746__13/HI _8841_/A sky130_fd_sc_hd__conb_1
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5040_ _5155_/B _5043_/A vssd1 vssd1 vccd1 vccd1 _5050_/C sky130_fd_sc_hd__or2_1
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6991_ _7347_/A _7347_/B _7347_/C _7347_/D vssd1 vssd1 vccd1 vccd1 _6991_/Y sky130_fd_sc_hd__nor4_1
XFILLER_53_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5942_ _5940_/Y _5941_/X _5953_/A vssd1 vssd1 vccd1 vccd1 _5955_/A sky130_fd_sc_hd__o21a_1
X_8730_ _8735_/CLK _8730_/D vssd1 vssd1 vccd1 vccd1 _8730_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_80_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5873_ _5873_/A vssd1 vssd1 vccd1 vccd1 _5981_/A sky130_fd_sc_hd__clkbuf_2
X_8661_ _8674_/CLK _8661_/D vssd1 vssd1 vccd1 vccd1 _8661_/Q sky130_fd_sc_hd__dfxtp_1
X_4824_ _4899_/A _4899_/B _4899_/C vssd1 vssd1 vccd1 vccd1 _4837_/B sky130_fd_sc_hd__nand3_2
XFILLER_61_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8592_ _8600_/CLK _8592_/D vssd1 vssd1 vccd1 vccd1 _8592_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7612_ _7613_/A _7613_/B _7613_/C vssd1 vssd1 vccd1 vccd1 _7614_/C sky130_fd_sc_hd__a21oi_1
X_7543_ _7543_/A _7543_/B vssd1 vssd1 vccd1 vccd1 _7543_/Y sky130_fd_sc_hd__nor2_1
X_4755_ _4755_/A vssd1 vssd1 vccd1 vccd1 _8614_/D sky130_fd_sc_hd__clkbuf_1
X_4686_ _4960_/A _5155_/A vssd1 vssd1 vccd1 vccd1 _4687_/B sky130_fd_sc_hd__nor2_1
X_7474_ _7509_/A _7505_/A _7496_/A vssd1 vssd1 vccd1 vccd1 _7491_/B sky130_fd_sc_hd__o21ai_1
X_6425_ _6425_/A _6425_/B vssd1 vssd1 vccd1 vccd1 _8681_/D sky130_fd_sc_hd__nor2_1
X_6356_ _6356_/A _6356_/B vssd1 vssd1 vccd1 vccd1 _6356_/Y sky130_fd_sc_hd__nor2_1
XFILLER_102_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5307_ _8637_/Q _5307_/B vssd1 vssd1 vccd1 vccd1 _5314_/C sky130_fd_sc_hd__and2_1
XFILLER_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6287_ _6186_/A _6186_/B _6286_/X vssd1 vssd1 vccd1 vccd1 _6288_/B sky130_fd_sc_hd__a21oi_1
X_8026_ _8026_/A _8026_/B vssd1 vssd1 vccd1 vccd1 _8031_/A sky130_fd_sc_hd__nand2_1
X_5238_ _5240_/B _5238_/B _5238_/C vssd1 vssd1 vccd1 vccd1 _5243_/B sky130_fd_sc_hd__or3_1
XFILLER_75_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5169_ _5169_/A _5245_/C vssd1 vssd1 vccd1 vccd1 _5170_/B sky130_fd_sc_hd__or2_1
XFILLER_84_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8830__97 vssd1 vssd1 vccd1 vccd1 _8830__97/HI _8654_/D sky130_fd_sc_hd__conb_1
XFILLER_71_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8928_ _8928_/A _4448_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[27] sky130_fd_sc_hd__ebufn_8
XFILLER_44_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8859_ _8859_/A _4367_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[28] sky130_fd_sc_hd__ebufn_8
XFILLER_71_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4540_ _4758_/A _4754_/B _4660_/B _4660_/A _5634_/B vssd1 vssd1 vccd1 vccd1 _4541_/D
+ sky130_fd_sc_hd__a2111o_1
X_4471_ _5453_/B vssd1 vssd1 vccd1 vccd1 _4720_/A sky130_fd_sc_hd__clkbuf_2
X_7190_ _7190_/A _7190_/B _7190_/C vssd1 vssd1 vccd1 vccd1 _7190_/X sky130_fd_sc_hd__or3_1
X_6210_ _6239_/A _6239_/B vssd1 vssd1 vccd1 vccd1 _6213_/A sky130_fd_sc_hd__xnor2_1
X_6141_ _6141_/A _6141_/B vssd1 vssd1 vccd1 vccd1 _6143_/C sky130_fd_sc_hd__nand2_1
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6072_ _6073_/A _6073_/B vssd1 vssd1 vccd1 vccd1 _6072_/X sky130_fd_sc_hd__or2_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5023_ _5028_/B _5015_/X _5017_/X _5022_/X vssd1 vssd1 vccd1 vccd1 _5023_/X sky130_fd_sc_hd__o211a_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6974_ _6973_/B _7366_/A _6973_/A vssd1 vssd1 vccd1 vccd1 _6975_/C sky130_fd_sc_hd__a21o_1
X_8713_ _8714_/CLK _8713_/D vssd1 vssd1 vccd1 vccd1 _8713_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5925_ _5925_/A _5925_/B vssd1 vssd1 vccd1 vccd1 _5926_/B sky130_fd_sc_hd__xnor2_1
X_8644_ _8681_/CLK _8644_/D vssd1 vssd1 vccd1 vccd1 _8644_/Q sky130_fd_sc_hd__dfxtp_1
X_5856_ _5856_/A _5856_/B vssd1 vssd1 vccd1 vccd1 _5856_/Y sky130_fd_sc_hd__nor2_1
X_4807_ _5220_/A vssd1 vssd1 vccd1 vccd1 _4916_/A sky130_fd_sc_hd__clkbuf_2
X_5787_ _6204_/B _5786_/Y _5893_/B vssd1 vssd1 vccd1 vccd1 _6211_/B sky130_fd_sc_hd__mux2_1
X_8575_ _8571_/A _7584_/X _8574_/Y _7544_/X vssd1 vssd1 vccd1 vccd1 _8734_/D sky130_fd_sc_hd__a211o_1
X_7526_ _7526_/A _7526_/B vssd1 vssd1 vccd1 vccd1 _7527_/B sky130_fd_sc_hd__and2_1
X_4738_ _6503_/A vssd1 vssd1 vccd1 vccd1 _7614_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_21_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7457_ _7457_/A _7457_/B vssd1 vssd1 vccd1 vccd1 _7458_/B sky130_fd_sc_hd__xnor2_1
X_4669_ _4763_/B vssd1 vssd1 vccd1 vccd1 _4752_/A sky130_fd_sc_hd__clkbuf_2
X_6408_ _8677_/Q _8676_/Q _8675_/Q vssd1 vssd1 vccd1 vccd1 _6413_/B sky130_fd_sc_hd__and3_1
XFILLER_79_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7388_ _7388_/A _7388_/B vssd1 vssd1 vccd1 vccd1 _7463_/B sky130_fd_sc_hd__xnor2_1
XFILLER_1_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6339_ _6339_/A vssd1 vssd1 vccd1 vccd1 _8668_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8009_ _8091_/A _8008_/Y _7985_/B _7921_/B vssd1 vssd1 vccd1 vccd1 _8020_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_29_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5710_ _5778_/A _5716_/A vssd1 vssd1 vccd1 vccd1 _5711_/B sky130_fd_sc_hd__xnor2_1
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6690_ _6690_/A vssd1 vssd1 vccd1 vccd1 _6876_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5641_ _5641_/A vssd1 vssd1 vccd1 vccd1 _5641_/Y sky130_fd_sc_hd__inv_2
X_8360_ _8351_/A _8351_/B _8359_/X vssd1 vssd1 vccd1 vccd1 _8437_/A sky130_fd_sc_hd__a21o_1
X_5572_ _5572_/A _5572_/B vssd1 vssd1 vccd1 vccd1 _5699_/B sky130_fd_sc_hd__xnor2_1
X_7311_ _6932_/A _6926_/A _7310_/X vssd1 vssd1 vccd1 vccd1 _7312_/B sky130_fd_sc_hd__o21ba_1
X_4523_ _5166_/A vssd1 vssd1 vccd1 vccd1 _4986_/B sky130_fd_sc_hd__clkbuf_2
X_8291_ _8291_/A _8291_/B vssd1 vssd1 vccd1 vccd1 _8292_/B sky130_fd_sc_hd__xor2_1
X_7242_ _7238_/A _7238_/B _7259_/A vssd1 vssd1 vccd1 vccd1 _7252_/A sky130_fd_sc_hd__a21bo_1
XFILLER_7_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4454_ _4455_/A vssd1 vssd1 vccd1 vccd1 _4454_/Y sky130_fd_sc_hd__inv_2
X_4385_ _4388_/A vssd1 vssd1 vccd1 vccd1 _4385_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7173_ _7173_/A _7173_/B vssd1 vssd1 vccd1 vccd1 _7175_/B sky130_fd_sc_hd__xor2_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6124_ _6133_/A _6124_/B vssd1 vssd1 vccd1 vccd1 _6126_/B sky130_fd_sc_hd__nand2_1
XFILLER_98_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6055_ _6051_/A _6055_/B vssd1 vssd1 vccd1 vccd1 _6089_/A sky130_fd_sc_hd__and2b_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5006_ _5016_/A _5121_/A vssd1 vssd1 vccd1 vccd1 _5007_/B sky130_fd_sc_hd__or2_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6957_ _6890_/A _6957_/B _7351_/A vssd1 vssd1 vccd1 vccd1 _6958_/C sky130_fd_sc_hd__and3b_1
XFILLER_81_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8800__67 vssd1 vssd1 vccd1 vccd1 _8800__67/HI _8909_/A sky130_fd_sc_hd__conb_1
XFILLER_81_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6888_ _6980_/A _7336_/S vssd1 vssd1 vccd1 vccd1 _6889_/B sky130_fd_sc_hd__xor2_1
X_5908_ _5933_/A _5933_/B vssd1 vssd1 vccd1 vccd1 _5926_/A sky130_fd_sc_hd__xor2_1
X_8627_ _8734_/CLK _8627_/D vssd1 vssd1 vccd1 vccd1 _8627_/Q sky130_fd_sc_hd__dfxtp_1
X_5839_ _5838_/A _5838_/C _5838_/B vssd1 vssd1 vccd1 vccd1 _5840_/B sky130_fd_sc_hd__o21ai_1
X_8558_ _8558_/A _8558_/B vssd1 vssd1 vccd1 vccd1 _8732_/D sky130_fd_sc_hd__nor2_1
X_7509_ _7509_/A _7509_/B vssd1 vssd1 vccd1 vccd1 _7510_/C sky130_fd_sc_hd__or2_1
X_8489_ _8489_/A _8489_/B vssd1 vssd1 vccd1 vccd1 _8490_/B sky130_fd_sc_hd__xnor2_1
XFILLER_5_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7860_ _7887_/A _7960_/B _7763_/B _7950_/B vssd1 vssd1 vccd1 vccd1 _7867_/A sky130_fd_sc_hd__a31o_1
XFILLER_35_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6811_ _6811_/A _6811_/B vssd1 vssd1 vccd1 vccd1 _6812_/B sky130_fd_sc_hd__nor2_1
XFILLER_63_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7791_ _8515_/C _8335_/A _7791_/C vssd1 vssd1 vccd1 vccd1 _7792_/B sky130_fd_sc_hd__nor3_1
X_6742_ _6742_/A _6742_/B vssd1 vssd1 vccd1 vccd1 _6742_/Y sky130_fd_sc_hd__nor2_1
XFILLER_50_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6673_ _6715_/A _6694_/B _6804_/A vssd1 vssd1 vccd1 vccd1 _6780_/A sky130_fd_sc_hd__nand3_1
X_5624_ _6039_/A _6037_/A vssd1 vssd1 vccd1 vccd1 _5676_/B sky130_fd_sc_hd__xnor2_1
X_8412_ _8412_/A _8412_/B vssd1 vssd1 vccd1 vccd1 _8414_/A sky130_fd_sc_hd__xnor2_1
X_8343_ _8343_/A _8343_/B vssd1 vssd1 vccd1 vccd1 _8345_/C sky130_fd_sc_hd__xnor2_1
X_5555_ _6134_/A _5896_/A _5556_/A _5554_/X vssd1 vssd1 vccd1 vccd1 _6024_/A sky130_fd_sc_hd__or4bb_1
X_4506_ _4787_/A _4749_/A _4786_/B _4786_/A vssd1 vssd1 vccd1 vccd1 _4511_/A sky130_fd_sc_hd__or4b_1
X_8274_ _8274_/A _8274_/B vssd1 vssd1 vccd1 vccd1 _8274_/Y sky130_fd_sc_hd__nor2_1
X_5486_ _8668_/Q vssd1 vssd1 vccd1 vccd1 _6338_/S sky130_fd_sc_hd__inv_2
X_4437_ _4437_/A vssd1 vssd1 vccd1 vccd1 _4437_/Y sky130_fd_sc_hd__inv_2
X_7225_ _7225_/A _7225_/B vssd1 vssd1 vccd1 vccd1 _7228_/B sky130_fd_sc_hd__xnor2_1
XFILLER_104_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7156_ _7156_/A _7156_/B vssd1 vssd1 vccd1 vccd1 _7159_/B sky130_fd_sc_hd__xnor2_1
X_4368_ _4369_/A vssd1 vssd1 vccd1 vccd1 _4368_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6107_ _5788_/A _6020_/Y _6071_/C _6071_/A vssd1 vssd1 vccd1 vccd1 _6108_/B sky130_fd_sc_hd__o22a_1
X_7087_ _7135_/A _7135_/B vssd1 vssd1 vccd1 vccd1 _7087_/X sky130_fd_sc_hd__or2_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6038_ _6038_/A _6066_/B vssd1 vssd1 vccd1 vccd1 _6039_/B sky130_fd_sc_hd__xnor2_1
XFILLER_26_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7989_ _8515_/A _7910_/A _8069_/A vssd1 vssd1 vccd1 vccd1 _7990_/A sky130_fd_sc_hd__mux2_1
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_2_0_wb_clk_i clkbuf_4_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _8600_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_45_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8791__58 vssd1 vssd1 vccd1 vccd1 _8791__58/HI _8900_/A sky130_fd_sc_hd__conb_1
XFILLER_32_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5340_ _5345_/C _5359_/A _5340_/C vssd1 vssd1 vccd1 vccd1 _5341_/A sky130_fd_sc_hd__and3b_1
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5271_ _5271_/A vssd1 vssd1 vccd1 vccd1 _5271_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_102_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7010_ _7010_/A _7010_/B _7063_/B vssd1 vssd1 vccd1 vccd1 _7314_/A sky130_fd_sc_hd__or3b_2
XFILLER_68_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7912_ _8008_/A _7912_/B vssd1 vssd1 vccd1 vccd1 _7985_/B sky130_fd_sc_hd__nor2_2
X_8892_ _8892_/A _4406_/Y vssd1 vssd1 vccd1 vccd1 io_out[29] sky130_fd_sc_hd__ebufn_8
XFILLER_36_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7843_ _7847_/A _7847_/B vssd1 vssd1 vccd1 vccd1 _7848_/A sky130_fd_sc_hd__nand2_1
X_4986_ _4986_/A _4986_/B _5073_/A _5231_/A vssd1 vssd1 vccd1 vccd1 _4987_/D sky130_fd_sc_hd__or4_1
XFILLER_63_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7774_ _7759_/A _7759_/B _7769_/X vssd1 vssd1 vccd1 vccd1 _7775_/B sky130_fd_sc_hd__a21oi_1
X_6725_ _6725_/A _6725_/B vssd1 vssd1 vccd1 vccd1 _6727_/A sky130_fd_sc_hd__xnor2_2
X_6656_ _6690_/A _6656_/B vssd1 vssd1 vccd1 vccd1 _6657_/A sky130_fd_sc_hd__and2b_1
XFILLER_31_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6587_ _6587_/A _7280_/C vssd1 vssd1 vccd1 vccd1 _6592_/A sky130_fd_sc_hd__xnor2_1
X_5607_ _5634_/A _7906_/B vssd1 vssd1 vccd1 vccd1 _5732_/A sky130_fd_sc_hd__nand2_1
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8326_ _8326_/A _8387_/A vssd1 vssd1 vccd1 vccd1 _8327_/B sky130_fd_sc_hd__xnor2_1
X_5538_ _5872_/A _5567_/B _5578_/A vssd1 vssd1 vccd1 vccd1 _5548_/A sky130_fd_sc_hd__and3_1
XFILLER_3_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8257_ _8257_/A _8257_/B vssd1 vssd1 vccd1 vccd1 _8259_/A sky130_fd_sc_hd__nor2_1
X_7208_ _7208_/A _7208_/B vssd1 vssd1 vccd1 vccd1 _7210_/B sky130_fd_sc_hd__xor2_1
X_5469_ _5470_/A _6598_/A vssd1 vssd1 vccd1 vccd1 _5493_/A sky130_fd_sc_hd__or2_1
XFILLER_59_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8188_ _8186_/Y _8183_/B _8187_/Y vssd1 vssd1 vccd1 vccd1 _8430_/A sky130_fd_sc_hd__a21oi_2
XFILLER_86_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7139_ _7181_/A _7181_/B _7139_/C vssd1 vssd1 vccd1 vccd1 _7141_/B sky130_fd_sc_hd__nand3_1
XFILLER_86_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4840_ _4990_/B _4849_/B vssd1 vssd1 vccd1 vccd1 _4999_/A sky130_fd_sc_hd__nor2_1
XFILLER_33_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6510_ _6565_/A _6511_/B vssd1 vssd1 vccd1 vccd1 _6510_/Y sky130_fd_sc_hd__nor2_1
XFILLER_60_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4771_ _7499_/A vssd1 vssd1 vccd1 vccd1 _4771_/X sky130_fd_sc_hd__buf_2
X_7490_ _7486_/Y _7394_/X _7489_/X vssd1 vssd1 vccd1 vccd1 _7491_/D sky130_fd_sc_hd__o21ba_1
X_6441_ _8687_/Q _6441_/B vssd1 vssd1 vccd1 vccd1 _6446_/C sky130_fd_sc_hd__and2_1
X_6372_ _6360_/A _6372_/B vssd1 vssd1 vccd1 vccd1 _6372_/X sky130_fd_sc_hd__and2b_1
X_5323_ _5323_/A vssd1 vssd1 vccd1 vccd1 _5323_/X sky130_fd_sc_hd__clkbuf_2
X_8111_ _8082_/A _8082_/B _8110_/Y vssd1 vssd1 vccd1 vccd1 _8190_/A sky130_fd_sc_hd__a21boi_2
X_5254_ _4718_/A _5080_/B _4715_/A _6746_/B vssd1 vssd1 vccd1 vccd1 _5255_/S sky130_fd_sc_hd__a22o_1
X_8042_ _8042_/A _8042_/B vssd1 vssd1 vccd1 vccd1 _8043_/B sky130_fd_sc_hd__xnor2_1
XFILLER_102_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5185_ _5185_/A _5185_/B _5227_/C _5185_/D vssd1 vssd1 vccd1 vccd1 _5186_/D sky130_fd_sc_hd__or4_1
XFILLER_83_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8875_ _8875_/A _4386_/Y vssd1 vssd1 vccd1 vccd1 io_out[12] sky130_fd_sc_hd__ebufn_8
XFILLER_83_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7826_ _7826_/A _7852_/A _7826_/C vssd1 vssd1 vccd1 vccd1 _7940_/A sky130_fd_sc_hd__or3_1
XFILLER_12_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4969_ _5130_/A _4969_/B vssd1 vssd1 vccd1 vccd1 _5139_/C sky130_fd_sc_hd__nand2_2
X_7757_ _7869_/A _7869_/B vssd1 vssd1 vccd1 vccd1 _7785_/A sky130_fd_sc_hd__xor2_1
X_6708_ _7254_/A _6999_/A vssd1 vssd1 vccd1 vccd1 _6708_/X sky130_fd_sc_hd__or2_1
X_7688_ _5453_/B _8732_/Q vssd1 vssd1 vccd1 vccd1 _7689_/B sky130_fd_sc_hd__and2b_1
X_6639_ _6639_/A _8621_/Q vssd1 vssd1 vccd1 vccd1 _6690_/A sky130_fd_sc_hd__and2_1
XFILLER_3_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8309_ _8309_/A _8367_/A vssd1 vssd1 vccd1 vccd1 _8310_/B sky130_fd_sc_hd__nand2_1
X_8736__3 vssd1 vssd1 vccd1 vccd1 _8736__3/HI _8831_/A sky130_fd_sc_hd__conb_1
XFILLER_93_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8761__28 vssd1 vssd1 vccd1 vccd1 _8761__28/HI _8856_/A sky130_fd_sc_hd__conb_1
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6990_ _6989_/A _6989_/B _6989_/C vssd1 vssd1 vccd1 vccd1 _7347_/D sky130_fd_sc_hd__a21oi_1
XFILLER_92_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5941_ _5941_/A _5941_/B _5941_/C vssd1 vssd1 vccd1 vccd1 _5941_/X sky130_fd_sc_hd__and3_1
XFILLER_25_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8660_ _8733_/CLK _8660_/D vssd1 vssd1 vccd1 vccd1 _8660_/Q sky130_fd_sc_hd__dfxtp_1
X_5872_ _5872_/A _5872_/B _5872_/C vssd1 vssd1 vccd1 vccd1 _5879_/A sky130_fd_sc_hd__and3_1
X_4823_ _4861_/B _4823_/B vssd1 vssd1 vccd1 vccd1 _4899_/C sky130_fd_sc_hd__xnor2_1
X_8591_ _8600_/CLK _8591_/D vssd1 vssd1 vccd1 vccd1 _8591_/Q sky130_fd_sc_hd__dfxtp_1
X_7611_ _7644_/A _7618_/B _7610_/X vssd1 vssd1 vccd1 vccd1 _7613_/C sky130_fd_sc_hd__a21oi_1
X_7542_ _7533_/A _7547_/S _7539_/Y _7546_/B _7548_/B vssd1 vssd1 vccd1 vccd1 _7543_/B
+ sky130_fd_sc_hd__a41o_1
X_4754_ _7550_/A _4754_/B _4754_/C vssd1 vssd1 vccd1 vccd1 _4755_/A sky130_fd_sc_hd__and3_1
X_7473_ _7473_/A _7473_/B vssd1 vssd1 vccd1 vccd1 _7496_/A sky130_fd_sc_hd__xnor2_1
X_4685_ _4914_/A vssd1 vssd1 vccd1 vccd1 _5155_/A sky130_fd_sc_hd__clkbuf_2
X_6424_ _6426_/A _6426_/C _6423_/X vssd1 vssd1 vccd1 vccd1 _6425_/B sky130_fd_sc_hd__o21ai_1
X_6355_ _6355_/A _6355_/B vssd1 vssd1 vccd1 vccd1 _6356_/B sky130_fd_sc_hd__nand2_1
X_5306_ _5306_/A vssd1 vssd1 vccd1 vccd1 _8636_/D sky130_fd_sc_hd__clkbuf_1
X_6286_ _6183_/B _6286_/B vssd1 vssd1 vccd1 vccd1 _6286_/X sky130_fd_sc_hd__and2b_1
XFILLER_102_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5237_ _5237_/A _5237_/B vssd1 vssd1 vccd1 vccd1 _5237_/Y sky130_fd_sc_hd__nor2_1
X_8025_ _8025_/A _8025_/B vssd1 vssd1 vccd1 vccd1 _8114_/A sky130_fd_sc_hd__nand2_1
XFILLER_102_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5168_ _4694_/A _5163_/X _5167_/X _5064_/A vssd1 vssd1 vccd1 vccd1 _5168_/X sky130_fd_sc_hd__a211o_1
XFILLER_83_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5099_ _5099_/A vssd1 vssd1 vccd1 vccd1 _5212_/A sky130_fd_sc_hd__clkbuf_2
X_8927_ _8927_/A _4447_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[26] sky130_fd_sc_hd__ebufn_8
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8858_ _8858_/A _4366_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[27] sky130_fd_sc_hd__ebufn_8
XFILLER_24_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7809_ _7813_/B _7809_/B vssd1 vssd1 vccd1 vccd1 _7901_/B sky130_fd_sc_hd__xnor2_1
XFILLER_12_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8806__73 vssd1 vssd1 vccd1 vccd1 _8806__73/HI _8915_/A sky130_fd_sc_hd__conb_1
XFILLER_58_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4470_ _8608_/Q vssd1 vssd1 vccd1 vccd1 _5453_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_7_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6140_ _6084_/A _6083_/B _6083_/C vssd1 vssd1 vccd1 vccd1 _6141_/B sky130_fd_sc_hd__o21ai_1
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6071_ _6071_/A _6204_/A _6071_/C vssd1 vssd1 vccd1 vccd1 _6073_/B sky130_fd_sc_hd__or3_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5022_ _5194_/C _5022_/B _5131_/A _5022_/D vssd1 vssd1 vccd1 vccd1 _5022_/X sky130_fd_sc_hd__or4_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6973_ _6973_/A _6973_/B _7366_/A vssd1 vssd1 vccd1 vccd1 _7366_/B sky130_fd_sc_hd__nand3_1
XFILLER_65_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8712_ _8714_/CLK _8712_/D vssd1 vssd1 vccd1 vccd1 _8712_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5924_ _5924_/A _5924_/B vssd1 vssd1 vccd1 vccd1 _5925_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8643_ _8710_/CLK _8643_/D vssd1 vssd1 vccd1 vccd1 _8643_/Q sky130_fd_sc_hd__dfxtp_1
X_5855_ _5848_/A _5848_/B _5854_/X vssd1 vssd1 vccd1 vccd1 _5930_/A sky130_fd_sc_hd__a21oi_1
X_4806_ _5226_/B vssd1 vssd1 vccd1 vccd1 _5220_/A sky130_fd_sc_hd__clkbuf_2
Xclkbuf_4_15_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8710_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_21_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5786_ _6204_/B _5997_/A vssd1 vssd1 vccd1 vccd1 _5786_/Y sky130_fd_sc_hd__nor2_1
X_8574_ _8574_/A _8574_/B vssd1 vssd1 vccd1 vccd1 _8574_/Y sky130_fd_sc_hd__nor2_1
X_7525_ _7526_/A _7532_/B vssd1 vssd1 vccd1 vccd1 _7535_/A sky130_fd_sc_hd__nor2_1
X_4737_ _4848_/C vssd1 vssd1 vccd1 vccd1 _4891_/A sky130_fd_sc_hd__clkbuf_2
X_7456_ _7456_/A _7456_/B vssd1 vssd1 vccd1 vccd1 _7457_/B sky130_fd_sc_hd__xnor2_1
X_4668_ _4668_/A _4668_/B _5028_/B _4698_/B vssd1 vssd1 vccd1 vccd1 _4763_/B sky130_fd_sc_hd__or4_1
X_6407_ _6407_/A vssd1 vssd1 vccd1 vccd1 _8676_/D sky130_fd_sc_hd__clkbuf_1
X_7387_ _7387_/A _7387_/B vssd1 vssd1 vccd1 vccd1 _7388_/B sky130_fd_sc_hd__nor2_1
X_4599_ _8585_/Q _4597_/A _4595_/X vssd1 vssd1 vccd1 vccd1 _4600_/B sky130_fd_sc_hd__o21ai_1
X_6338_ _5397_/A _5398_/A _6338_/S vssd1 vssd1 vccd1 vccd1 _6339_/A sky130_fd_sc_hd__mux2_1
X_6269_ _6178_/A _6178_/B _6268_/X vssd1 vssd1 vccd1 vccd1 _6276_/A sky130_fd_sc_hd__a21oi_1
XFILLER_57_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8008_ _8008_/A _8008_/B vssd1 vssd1 vccd1 vccd1 _8008_/Y sky130_fd_sc_hd__nor2_1
XFILLER_84_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5640_ _5742_/A _5859_/A vssd1 vssd1 vccd1 vccd1 _5640_/Y sky130_fd_sc_hd__nand2_1
X_5571_ _5571_/A _5571_/B vssd1 vssd1 vccd1 vccd1 _5572_/B sky130_fd_sc_hd__xor2_1
X_7310_ _7310_/A _7336_/S _7369_/B vssd1 vssd1 vccd1 vccd1 _7310_/X sky130_fd_sc_hd__and3_1
X_4522_ _4522_/A vssd1 vssd1 vccd1 vccd1 _5166_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_8290_ _8290_/A _8362_/B vssd1 vssd1 vccd1 vccd1 _8292_/A sky130_fd_sc_hd__xnor2_1
X_4453_ _4455_/A vssd1 vssd1 vccd1 vccd1 _4453_/Y sky130_fd_sc_hd__inv_2
X_7241_ _7258_/A _7258_/B vssd1 vssd1 vccd1 vccd1 _7259_/A sky130_fd_sc_hd__or2_1
X_4384_ _4388_/A vssd1 vssd1 vccd1 vccd1 _4384_/Y sky130_fd_sc_hd__inv_2
X_7172_ _7454_/A _7172_/B _7172_/C vssd1 vssd1 vccd1 vccd1 _7234_/A sky130_fd_sc_hd__and3_1
XFILLER_98_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6123_ _6316_/B _6098_/S _5947_/X _6121_/Y _6122_/X vssd1 vssd1 vccd1 vccd1 _6124_/B
+ sky130_fd_sc_hd__a32o_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6054_ _6056_/B _6056_/A vssd1 vssd1 vccd1 vccd1 _6091_/A sky130_fd_sc_hd__and2b_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5005_ _5166_/A _5215_/B _5155_/C _5003_/X _5120_/D vssd1 vssd1 vccd1 vccd1 _5005_/X
+ sky130_fd_sc_hd__o32a_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8797__64 vssd1 vssd1 vccd1 vccd1 _8797__64/HI _8906_/A sky130_fd_sc_hd__conb_1
XFILLER_38_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6956_ _6890_/A _7350_/B _7352_/C _6876_/B vssd1 vssd1 vccd1 vccd1 _6958_/B sky130_fd_sc_hd__o22a_1
XFILLER_41_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5907_ _5907_/A _5907_/B vssd1 vssd1 vccd1 vccd1 _5933_/B sky130_fd_sc_hd__xnor2_2
XFILLER_22_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6887_ _7000_/B vssd1 vssd1 vccd1 vccd1 _7336_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_34_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8626_ _8734_/CLK _8626_/D vssd1 vssd1 vccd1 vccd1 _8626_/Q sky130_fd_sc_hd__dfxtp_1
X_5838_ _5838_/A _5838_/B _5838_/C vssd1 vssd1 vccd1 vccd1 _5838_/Y sky130_fd_sc_hd__nor3_1
X_8557_ _8556_/Y _8553_/A _8578_/A vssd1 vssd1 vccd1 vccd1 _8558_/B sky130_fd_sc_hd__mux2_1
X_5769_ _5769_/A _5850_/B vssd1 vssd1 vccd1 vccd1 _6018_/B sky130_fd_sc_hd__xnor2_1
X_7508_ _7509_/A _7509_/B vssd1 vssd1 vccd1 vccd1 _7510_/B sky130_fd_sc_hd__nand2_1
XFILLER_5_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8488_ _8422_/A _8422_/B _8487_/X vssd1 vssd1 vccd1 vccd1 _8490_/A sky130_fd_sc_hd__a21oi_1
X_7439_ _7439_/A _7439_/B vssd1 vssd1 vccd1 vccd1 _7439_/Y sky130_fd_sc_hd__nor2_1
XFILLER_30_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6810_ _6826_/A vssd1 vssd1 vccd1 vccd1 _6811_/A sky130_fd_sc_hd__inv_2
XFILLER_63_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7790_ _8203_/B _8331_/A vssd1 vssd1 vccd1 vccd1 _7791_/C sky130_fd_sc_hd__nor2_1
X_6741_ _6742_/A _6742_/B vssd1 vssd1 vccd1 vccd1 _7091_/B sky130_fd_sc_hd__xor2_1
X_6672_ _6672_/A vssd1 vssd1 vccd1 vccd1 _6804_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5623_ _5952_/A _5967_/A vssd1 vssd1 vccd1 vccd1 _6037_/A sky130_fd_sc_hd__nor2_1
X_8411_ _7963_/X _8410_/Y _8411_/S vssd1 vssd1 vccd1 vccd1 _8412_/B sky130_fd_sc_hd__mux2_1
X_8342_ _8342_/A _8342_/B vssd1 vssd1 vccd1 vccd1 _8343_/B sky130_fd_sc_hd__nor2_1
X_5554_ _5557_/B _5552_/C _5552_/A vssd1 vssd1 vccd1 vccd1 _5554_/X sky130_fd_sc_hd__a21o_1
X_4505_ _4660_/A vssd1 vssd1 vccd1 vccd1 _4786_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_8273_ _8257_/B _8259_/B _8257_/A vssd1 vssd1 vccd1 vccd1 _8353_/A sky130_fd_sc_hd__o21ba_1
X_5485_ _5780_/A _5874_/B vssd1 vssd1 vccd1 vccd1 _5498_/A sky130_fd_sc_hd__nand2_1
X_4436_ _4437_/A vssd1 vssd1 vccd1 vccd1 _4436_/Y sky130_fd_sc_hd__inv_2
X_7224_ _7223_/A _7245_/A vssd1 vssd1 vccd1 vccd1 _7228_/A sky130_fd_sc_hd__and2b_1
XFILLER_6_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4367_ _4369_/A vssd1 vssd1 vccd1 vccd1 _4367_/Y sky130_fd_sc_hd__inv_2
X_7155_ _7190_/B _7190_/C _7190_/A vssd1 vssd1 vccd1 vccd1 _7159_/A sky130_fd_sc_hd__o21ba_1
XFILLER_98_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6106_ _6106_/A _6106_/B vssd1 vssd1 vccd1 vccd1 _6116_/A sky130_fd_sc_hd__or2_1
XFILLER_98_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7086_ _7169_/A _7348_/B _7170_/A vssd1 vssd1 vccd1 vccd1 _7135_/B sky130_fd_sc_hd__and3_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6037_ _6037_/A _6037_/B vssd1 vssd1 vccd1 vccd1 _6066_/B sky130_fd_sc_hd__xnor2_1
XFILLER_39_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7988_ _7988_/A _8146_/B vssd1 vssd1 vccd1 vccd1 _8069_/A sky130_fd_sc_hd__nand2_2
XFILLER_26_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6939_ _7039_/A _6939_/B vssd1 vssd1 vccd1 vccd1 _7046_/A sky130_fd_sc_hd__xnor2_1
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8609_ _8733_/CLK _8609_/D vssd1 vssd1 vccd1 vccd1 _8609_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5270_ _8725_/Q _5258_/X _5269_/X _5267_/X vssd1 vssd1 vccd1 vccd1 _8626_/D sky130_fd_sc_hd__o211a_1
XFILLER_99_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7911_ _7798_/B _8065_/B _8243_/B vssd1 vssd1 vccd1 vccd1 _7912_/B sky130_fd_sc_hd__a21oi_1
X_8891_ _8891_/A _4405_/Y vssd1 vssd1 vccd1 vccd1 io_out[28] sky130_fd_sc_hd__ebufn_8
X_8767__34 vssd1 vssd1 vccd1 vccd1 _8767__34/HI _8862_/A sky130_fd_sc_hd__conb_1
XFILLER_83_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7842_ _8514_/A _8514_/B _8518_/B vssd1 vssd1 vccd1 vccd1 _7847_/B sky130_fd_sc_hd__and3_1
X_4985_ _5009_/B _5172_/B _4987_/C _4984_/X vssd1 vssd1 vccd1 vccd1 _4985_/X sky130_fd_sc_hd__o31a_1
XFILLER_51_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7773_ _7773_/A _7955_/C _7955_/D vssd1 vssd1 vccd1 vccd1 _7972_/A sky130_fd_sc_hd__or3_2
X_6724_ _6724_/A _6724_/B vssd1 vssd1 vccd1 vccd1 _6725_/B sky130_fd_sc_hd__xnor2_2
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6655_ _6655_/A vssd1 vssd1 vccd1 vccd1 _6715_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6586_ _7275_/A _6893_/B _6586_/C vssd1 vssd1 vccd1 vccd1 _7280_/C sky130_fd_sc_hd__and3_1
X_5606_ _5940_/B _6028_/B vssd1 vssd1 vccd1 vccd1 _5682_/A sky130_fd_sc_hd__nor2_2
X_8325_ _8325_/A _8325_/B vssd1 vssd1 vccd1 vccd1 _8387_/A sky130_fd_sc_hd__xnor2_1
X_5537_ _5874_/B _5780_/B _5780_/C vssd1 vssd1 vccd1 vccd1 _5578_/A sky130_fd_sc_hd__and3_1
XFILLER_11_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8256_ _8256_/A _8256_/B _8256_/C vssd1 vssd1 vccd1 vccd1 _8257_/B sky130_fd_sc_hd__nor3_1
XFILLER_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7207_ _7234_/A _7234_/B _7235_/B vssd1 vssd1 vccd1 vccd1 _7210_/A sky130_fd_sc_hd__or3_1
X_5468_ _8610_/Q vssd1 vssd1 vccd1 vccd1 _6598_/A sky130_fd_sc_hd__buf_2
X_8187_ _8187_/A _8187_/B vssd1 vssd1 vccd1 vccd1 _8187_/Y sky130_fd_sc_hd__nor2_1
X_5399_ _8656_/Q _5400_/A vssd1 vssd1 vccd1 vccd1 _5401_/A sky130_fd_sc_hd__or2b_1
X_4419_ _4419_/A vssd1 vssd1 vccd1 vccd1 _4419_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7138_ _7145_/B _7138_/B vssd1 vssd1 vccd1 vccd1 _7139_/C sky130_fd_sc_hd__xor2_1
XFILLER_100_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7069_ _7069_/A _7211_/A _7068_/X vssd1 vssd1 vccd1 vccd1 _7167_/A sky130_fd_sc_hd__nor3b_1
XFILLER_100_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4770_ _4808_/A vssd1 vssd1 vccd1 vccd1 _4774_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6440_ _6440_/A vssd1 vssd1 vccd1 vccd1 _8686_/D sky130_fd_sc_hd__clkbuf_1
X_6371_ _5398_/X _6370_/Y _8673_/Q _4582_/B vssd1 vssd1 vccd1 vccd1 _8673_/D sky130_fd_sc_hd__o2bb2a_1
X_5322_ _8641_/Q _8640_/Q _5322_/C vssd1 vssd1 vccd1 vccd1 _5328_/C sky130_fd_sc_hd__and3_1
X_8110_ _8110_/A _8110_/B vssd1 vssd1 vccd1 vccd1 _8110_/Y sky130_fd_sc_hd__nand2_1
X_5253_ _5149_/S _5158_/X _5191_/X _5252_/X vssd1 vssd1 vccd1 vccd1 _5253_/X sky130_fd_sc_hd__a31o_1
X_8041_ _8041_/A _8041_/B vssd1 vssd1 vccd1 vccd1 _8042_/B sky130_fd_sc_hd__xnor2_1
X_5184_ _4906_/A _4904_/A _4937_/A vssd1 vssd1 vccd1 vccd1 _5185_/D sky130_fd_sc_hd__a21oi_1
XFILLER_3_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8874_ _8874_/A _4385_/Y vssd1 vssd1 vccd1 vccd1 io_out[11] sky130_fd_sc_hd__ebufn_8
XFILLER_83_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7825_ _7825_/A _7825_/B vssd1 vssd1 vccd1 vccd1 _7826_/C sky130_fd_sc_hd__and2_1
XFILLER_12_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4968_ _5244_/A vssd1 vssd1 vccd1 vccd1 _5130_/A sky130_fd_sc_hd__buf_2
X_7756_ _7759_/A _7759_/B _7769_/A vssd1 vssd1 vccd1 vccd1 _7869_/B sky130_fd_sc_hd__a21oi_4
XFILLER_51_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6707_ _6800_/A vssd1 vssd1 vccd1 vccd1 _7409_/A sky130_fd_sc_hd__clkbuf_2
X_4899_ _4899_/A _4899_/B _4899_/C vssd1 vssd1 vccd1 vccd1 _5087_/B sky130_fd_sc_hd__and3_1
X_7687_ _8732_/Q _8608_/Q vssd1 vssd1 vccd1 vccd1 _7689_/A sky130_fd_sc_hd__and2b_2
X_6638_ _6659_/A _6652_/B _6652_/C _6637_/Y vssd1 vssd1 vccd1 vccd1 _6689_/A sky130_fd_sc_hd__a31o_2
X_6569_ _6588_/A _6578_/B vssd1 vssd1 vccd1 vccd1 _6699_/A sky130_fd_sc_hd__xor2_1
X_8308_ _8308_/A _8309_/A vssd1 vssd1 vccd1 vccd1 _8312_/B sky130_fd_sc_hd__or2_1
XFILLER_78_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8239_ _8239_/A _8300_/B vssd1 vssd1 vccd1 vccd1 _8240_/B sky130_fd_sc_hd__xnor2_1
XFILLER_78_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5940_ _6120_/A _5940_/B vssd1 vssd1 vccd1 vccd1 _5940_/Y sky130_fd_sc_hd__nor2_1
XFILLER_80_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5871_ _5808_/A _5808_/B _5870_/X vssd1 vssd1 vccd1 vccd1 _5906_/A sky130_fd_sc_hd__a21oi_2
XFILLER_33_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7610_ _7644_/A _7618_/B _7604_/X vssd1 vssd1 vccd1 vccd1 _7610_/X sky130_fd_sc_hd__o21a_1
X_4822_ _4822_/A _4822_/B vssd1 vssd1 vccd1 vccd1 _4899_/A sky130_fd_sc_hd__or2_1
X_8590_ _8600_/CLK _8590_/D vssd1 vssd1 vccd1 vccd1 _8590_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7541_ _7533_/A _7547_/S _7539_/Y _7546_/B vssd1 vssd1 vccd1 vccd1 _7543_/A sky130_fd_sc_hd__a22oi_1
X_4753_ _4758_/B _4752_/X _4749_/A _5265_/A vssd1 vssd1 vccd1 vccd1 _4754_/C sky130_fd_sc_hd__a2bb2o_1
X_7472_ _7472_/A _7266_/X vssd1 vssd1 vccd1 vccd1 _7473_/A sky130_fd_sc_hd__or2b_1
X_6423_ _6464_/B vssd1 vssd1 vccd1 vccd1 _6423_/X sky130_fd_sc_hd__buf_4
X_4684_ _5175_/A vssd1 vssd1 vccd1 vccd1 _4914_/A sky130_fd_sc_hd__clkbuf_2
X_6354_ _6354_/A _6354_/B vssd1 vssd1 vccd1 vccd1 _6356_/A sky130_fd_sc_hd__nand2_1
X_5305_ _5307_/B _5359_/A _5305_/C vssd1 vssd1 vccd1 vccd1 _5306_/A sky130_fd_sc_hd__and3b_1
X_6285_ _6181_/A _6181_/B _6182_/B _6182_/A vssd1 vssd1 vccd1 vccd1 _6288_/A sky130_fd_sc_hd__a2bb2o_1
X_5236_ _8603_/Q _5245_/C _5236_/C _5245_/D vssd1 vssd1 vccd1 vccd1 _5236_/X sky130_fd_sc_hd__or4_1
X_8024_ _8024_/A _8024_/B vssd1 vssd1 vccd1 vccd1 _8112_/B sky130_fd_sc_hd__nand2_2
XFILLER_84_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5167_ _5096_/B _5165_/X _5166_/X _5107_/C _5053_/A vssd1 vssd1 vccd1 vccd1 _5167_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_68_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5098_ _5223_/B _5109_/B vssd1 vssd1 vccd1 vccd1 _5139_/D sky130_fd_sc_hd__or2_1
XFILLER_83_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8926_ _8926_/A _4446_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[25] sky130_fd_sc_hd__ebufn_8
XFILLER_71_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8857_ _8857_/A _4365_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[26] sky130_fd_sc_hd__ebufn_8
XFILLER_52_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7808_ _7818_/A _7903_/C vssd1 vssd1 vccd1 vccd1 _7809_/B sky130_fd_sc_hd__xnor2_1
X_7739_ _7739_/A _7738_/X vssd1 vssd1 vccd1 vccd1 _7742_/A sky130_fd_sc_hd__or2b_1
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8821__88 vssd1 vssd1 vccd1 vccd1 _8821__88/HI _8930_/A sky130_fd_sc_hd__conb_1
XFILLER_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6070_ _6118_/A _6070_/B vssd1 vssd1 vccd1 vccd1 _6071_/C sky130_fd_sc_hd__or2_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5021_ _5038_/A _5062_/C _5179_/B _5009_/B vssd1 vssd1 vccd1 vccd1 _5022_/D sky130_fd_sc_hd__o31a_1
XFILLER_66_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8711_ _8715_/CLK _8711_/D vssd1 vssd1 vccd1 vccd1 _8711_/Q sky130_fd_sc_hd__dfxtp_1
X_6972_ _7352_/A _7350_/A _6972_/C vssd1 vssd1 vccd1 vccd1 _7366_/A sky130_fd_sc_hd__or3_1
XFILLER_19_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5923_ _5923_/A _5923_/B vssd1 vssd1 vccd1 vccd1 _5925_/A sky130_fd_sc_hd__nor2_1
X_8642_ _8681_/CLK _8642_/D vssd1 vssd1 vccd1 vccd1 _8642_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5854_ _5830_/A _5854_/B vssd1 vssd1 vccd1 vccd1 _5854_/X sky130_fd_sc_hd__and2b_1
XFILLER_21_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4805_ _4765_/A _4790_/Y _4799_/X _4803_/X _4804_/X vssd1 vssd1 vccd1 vccd1 _4805_/X
+ sky130_fd_sc_hd__o2111a_1
X_8573_ _8573_/A _8573_/B vssd1 vssd1 vccd1 vccd1 _8574_/B sky130_fd_sc_hd__xnor2_1
X_7524_ _7520_/A _5308_/X _6508_/X _7523_/X vssd1 vssd1 vccd1 vccd1 _8711_/D sky130_fd_sc_hd__a22o_1
X_5785_ _5992_/B vssd1 vssd1 vccd1 vccd1 _5997_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4736_ _8612_/Q vssd1 vssd1 vccd1 vccd1 _4848_/C sky130_fd_sc_hd__inv_2
X_7455_ _7355_/B _7455_/B vssd1 vssd1 vccd1 vccd1 _7456_/B sky130_fd_sc_hd__and2b_1
X_4667_ _5079_/A _5205_/A vssd1 vssd1 vccd1 vccd1 _4698_/B sky130_fd_sc_hd__nand2_2
X_7386_ _7429_/B _7385_/B _7385_/C vssd1 vssd1 vccd1 vccd1 _7387_/B sky130_fd_sc_hd__o21a_1
X_6406_ _6397_/A _6406_/B _6406_/C vssd1 vssd1 vccd1 vccd1 _6407_/A sky130_fd_sc_hd__and3b_1
XFILLER_1_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6337_ _6324_/X _6336_/X _6325_/X _8667_/Q vssd1 vssd1 vccd1 vccd1 _8667_/D sky130_fd_sc_hd__o2bb2a_1
X_4598_ _8584_/Q _8585_/Q _4598_/C vssd1 vssd1 vccd1 vccd1 _4604_/C sky130_fd_sc_hd__and3_1
X_6268_ _6177_/A _6268_/B vssd1 vssd1 vccd1 vccd1 _6268_/X sky130_fd_sc_hd__and2b_1
XFILLER_88_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5219_ _5120_/B _5212_/X _4914_/A vssd1 vssd1 vccd1 vccd1 _5220_/D sky130_fd_sc_hd__o21a_1
XFILLER_69_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6199_ _6199_/A _6006_/A vssd1 vssd1 vccd1 vccd1 _6201_/A sky130_fd_sc_hd__or2b_1
X_8007_ _8008_/A _8008_/B vssd1 vssd1 vccd1 vccd1 _8091_/A sky130_fd_sc_hd__and2_1
XFILLER_29_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8909_ _8909_/A _4418_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[8] sky130_fd_sc_hd__ebufn_8
XFILLER_40_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5570_ _6204_/A _5781_/A _5569_/X vssd1 vssd1 vccd1 vccd1 _5571_/B sky130_fd_sc_hd__a21oi_1
X_4521_ _5171_/A _5199_/A vssd1 vssd1 vccd1 vccd1 _4522_/A sky130_fd_sc_hd__or2_1
X_4452_ _4455_/A vssd1 vssd1 vccd1 vccd1 _4452_/Y sky130_fd_sc_hd__inv_2
X_7240_ _7280_/B _7069_/A _7239_/X vssd1 vssd1 vccd1 vccd1 _7258_/B sky130_fd_sc_hd__a21o_1
XFILLER_104_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4383_ _4401_/A vssd1 vssd1 vccd1 vccd1 _4388_/A sky130_fd_sc_hd__buf_4
X_7171_ _7275_/A _7213_/B _7213_/D vssd1 vssd1 vccd1 vccd1 _7182_/A sky130_fd_sc_hd__or3b_1
XFILLER_98_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6122_ _6122_/A _6122_/B vssd1 vssd1 vccd1 vccd1 _6122_/X sky130_fd_sc_hd__or2_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6053_ _6085_/A _6085_/B _6052_/X vssd1 vssd1 vccd1 vccd1 _6056_/A sky130_fd_sc_hd__a21o_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5004_ _5171_/A _5243_/A vssd1 vssd1 vccd1 vccd1 _5120_/D sky130_fd_sc_hd__nand2_2
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6955_ _7172_/B _7083_/B vssd1 vssd1 vccd1 vccd1 _7348_/C sky130_fd_sc_hd__and2_1
XFILLER_81_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5906_ _5906_/A _5965_/B vssd1 vssd1 vccd1 vccd1 _5907_/B sky130_fd_sc_hd__xnor2_2
X_6886_ _6730_/A _6730_/B _6813_/A _7332_/A vssd1 vssd1 vccd1 vccd1 _7000_/B sky130_fd_sc_hd__a211o_1
X_8625_ _8734_/CLK _8625_/D vssd1 vssd1 vccd1 vccd1 _8625_/Q sky130_fd_sc_hd__dfxtp_1
X_5837_ _6194_/A _5837_/B vssd1 vssd1 vccd1 vccd1 _5838_/C sky130_fd_sc_hd__nor2_1
XFILLER_22_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8556_ _8556_/A _8562_/B vssd1 vssd1 vccd1 vccd1 _8556_/Y sky130_fd_sc_hd__xnor2_1
X_5768_ _5847_/A _5768_/B vssd1 vssd1 vccd1 vccd1 _5850_/B sky130_fd_sc_hd__nand2_1
X_4719_ _4719_/A _5034_/B vssd1 vssd1 vccd1 vccd1 _4726_/B sky130_fd_sc_hd__nor2_1
X_7507_ _7499_/X _8707_/Q _7497_/X _7506_/X vssd1 vssd1 vccd1 vccd1 _8707_/D sky130_fd_sc_hd__o22a_1
X_8487_ _8423_/A _8487_/B vssd1 vssd1 vccd1 vccd1 _8487_/X sky130_fd_sc_hd__and2b_1
X_7438_ _7439_/A _7439_/B vssd1 vssd1 vccd1 vccd1 _7438_/Y sky130_fd_sc_hd__nand2_1
X_5699_ _5699_/A _5699_/B vssd1 vssd1 vccd1 vccd1 _5699_/Y sky130_fd_sc_hd__nand2_1
X_7369_ _7369_/A _7369_/B vssd1 vssd1 vccd1 vccd1 _7372_/A sky130_fd_sc_hd__nor2_1
XFILLER_89_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6740_ _6793_/C _7127_/A vssd1 vssd1 vccd1 vccd1 _6742_/B sky130_fd_sc_hd__xnor2_1
XFILLER_63_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6671_ _7074_/B _6734_/B _7074_/C _7130_/A vssd1 vssd1 vccd1 vccd1 _6672_/A sky130_fd_sc_hd__or4b_2
X_5622_ _5630_/A _5630_/B vssd1 vssd1 vccd1 vccd1 _5967_/A sky130_fd_sc_hd__xor2_4
X_8410_ _8410_/A _8410_/B vssd1 vssd1 vccd1 vccd1 _8410_/Y sky130_fd_sc_hd__nor2_1
X_5553_ _6070_/B vssd1 vssd1 vccd1 vccd1 _6134_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_8341_ _8415_/A _8341_/B _8413_/B vssd1 vssd1 vccd1 vccd1 _8342_/B sky130_fd_sc_hd__and3_1
X_4504_ _7737_/B vssd1 vssd1 vccd1 vccd1 _4660_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_8272_ _8262_/A _8262_/B _8271_/Y vssd1 vssd1 vccd1 vccd1 _8431_/A sky130_fd_sc_hd__a21o_1
X_5484_ _5892_/A _5513_/B vssd1 vssd1 vccd1 vccd1 _5500_/A sky130_fd_sc_hd__xnor2_1
X_4435_ _4437_/A vssd1 vssd1 vccd1 vccd1 _4435_/Y sky130_fd_sc_hd__inv_2
X_7223_ _7223_/A _7223_/B _7223_/C vssd1 vssd1 vccd1 vccd1 _7245_/A sky130_fd_sc_hd__or3_1
X_4366_ _4369_/A vssd1 vssd1 vccd1 vccd1 _4366_/Y sky130_fd_sc_hd__inv_2
X_7154_ _7185_/A _7154_/B _7154_/C vssd1 vssd1 vccd1 vccd1 _7190_/A sky130_fd_sc_hd__and3b_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6105_ _6316_/B _5682_/A _5940_/Y _6101_/A _6102_/X vssd1 vssd1 vccd1 vccd1 _6106_/B
+ sky130_fd_sc_hd__a2111oi_1
XFILLER_100_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7085_ _7172_/C _7085_/B vssd1 vssd1 vccd1 vccd1 _7135_/A sky130_fd_sc_hd__xor2_1
XFILLER_58_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6036_ _6036_/A _6036_/B vssd1 vssd1 vccd1 vccd1 _6063_/A sky130_fd_sc_hd__xnor2_1
XFILLER_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7987_ _7802_/B _7804_/B _7906_/X vssd1 vssd1 vccd1 vccd1 _8146_/B sky130_fd_sc_hd__a21oi_4
XFILLER_26_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6938_ _7023_/B _6938_/B vssd1 vssd1 vccd1 vccd1 _6939_/B sky130_fd_sc_hd__xnor2_1
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6869_ _6869_/A _6869_/B vssd1 vssd1 vccd1 vccd1 _6901_/B sky130_fd_sc_hd__nand2_1
X_8608_ _8733_/CLK _8608_/D vssd1 vssd1 vccd1 vccd1 _8608_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8539_ _8716_/Q _8540_/A vssd1 vssd1 vccd1 vccd1 _8541_/A sky130_fd_sc_hd__or2b_1
XFILLER_41_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8890_ _8890_/A _4404_/Y vssd1 vssd1 vccd1 vccd1 io_out[27] sky130_fd_sc_hd__ebufn_8
XFILLER_83_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7910_ _7910_/A vssd1 vssd1 vccd1 vccd1 _8243_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7841_ _7841_/A _7841_/B vssd1 vssd1 vccd1 vccd1 _8518_/B sky130_fd_sc_hd__xor2_1
XFILLER_23_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8782__49 vssd1 vssd1 vccd1 vccd1 _8782__49/HI _8891_/A sky130_fd_sc_hd__conb_1
X_4984_ _5175_/C _5188_/C _4984_/C _4984_/D vssd1 vssd1 vccd1 vccd1 _4984_/X sky130_fd_sc_hd__or4_1
X_7772_ _7771_/A _7771_/C _7771_/B vssd1 vssd1 vccd1 vccd1 _7955_/D sky130_fd_sc_hd__a21oi_1
X_6723_ _6774_/S _6780_/B _6722_/X vssd1 vssd1 vccd1 vccd1 _6724_/B sky130_fd_sc_hd__a21o_1
XFILLER_23_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6654_ _6870_/A _6870_/B vssd1 vssd1 vccd1 vccd1 _6655_/A sky130_fd_sc_hd__and2_1
X_5605_ _5605_/A _5605_/B vssd1 vssd1 vccd1 vccd1 _6028_/B sky130_fd_sc_hd__xor2_4
X_6585_ _6578_/B _7430_/A _7128_/A vssd1 vssd1 vccd1 vccd1 _6586_/C sky130_fd_sc_hd__o21ai_1
XFILLER_11_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5536_ _5558_/B _5535_/C _5535_/A vssd1 vssd1 vccd1 vccd1 _5550_/B sky130_fd_sc_hd__a21oi_1
X_8324_ _8324_/A _8324_/B vssd1 vssd1 vccd1 vccd1 _8325_/B sky130_fd_sc_hd__nor2_1
X_8255_ _8256_/A _8256_/B _8256_/C vssd1 vssd1 vccd1 vccd1 _8257_/A sky130_fd_sc_hd__o21a_1
X_5467_ _8673_/Q vssd1 vssd1 vccd1 vccd1 _5470_/A sky130_fd_sc_hd__inv_2
X_7206_ _7213_/D _7206_/B vssd1 vssd1 vccd1 vccd1 _7235_/B sky130_fd_sc_hd__xnor2_1
X_4418_ _4419_/A vssd1 vssd1 vccd1 vccd1 _4418_/Y sky130_fd_sc_hd__inv_2
X_8186_ _8186_/A vssd1 vssd1 vccd1 vccd1 _8186_/Y sky130_fd_sc_hd__inv_2
X_5398_ _5398_/A vssd1 vssd1 vccd1 vccd1 _5398_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_98_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7137_ _7128_/A _7352_/B _6880_/X _7169_/A vssd1 vssd1 vccd1 vccd1 _7181_/B sky130_fd_sc_hd__o211a_1
X_4349_ _4351_/A vssd1 vssd1 vccd1 vccd1 _4349_/Y sky130_fd_sc_hd__inv_2
X_7068_ _7068_/A _7270_/A vssd1 vssd1 vccd1 vccd1 _7068_/X sky130_fd_sc_hd__xor2_1
XFILLER_86_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6019_ _6019_/A _6019_/B vssd1 vssd1 vccd1 vccd1 _6069_/A sky130_fd_sc_hd__xnor2_1
XFILLER_46_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6370_ _6370_/A _6370_/B vssd1 vssd1 vccd1 vccd1 _6370_/Y sky130_fd_sc_hd__xnor2_1
X_5321_ _5321_/A _5321_/B vssd1 vssd1 vccd1 vccd1 _8640_/D sky130_fd_sc_hd__nor2_1
XFILLER_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8040_ _8040_/A _8040_/B vssd1 vssd1 vccd1 vccd1 _8041_/B sky130_fd_sc_hd__nor2_1
X_5252_ _5096_/B _5251_/X _5149_/S vssd1 vssd1 vccd1 vccd1 _5252_/X sky130_fd_sc_hd__o21ba_1
X_8827__94 vssd1 vssd1 vccd1 vccd1 _8827__94/HI _8936_/A sky130_fd_sc_hd__conb_1
X_5183_ _5199_/A _5240_/B _5183_/C _5244_/C vssd1 vssd1 vccd1 vccd1 _5183_/X sky130_fd_sc_hd__or4_1
XFILLER_68_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8873_ _8873_/A _4384_/Y vssd1 vssd1 vccd1 vccd1 io_out[10] sky130_fd_sc_hd__ebufn_8
XFILLER_71_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7824_ _7825_/A _7825_/B vssd1 vssd1 vccd1 vccd1 _7852_/A sky130_fd_sc_hd__nor2_1
X_4967_ _5223_/D _5188_/C _5180_/D _5172_/A _5214_/A vssd1 vssd1 vccd1 vccd1 _4970_/C
+ sky130_fd_sc_hd__o32a_1
X_7755_ _7775_/A _7769_/B vssd1 vssd1 vccd1 vccd1 _7869_/A sky130_fd_sc_hd__or2_2
XFILLER_51_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6706_ _7099_/A _7099_/B _7099_/C _6651_/B _7103_/A vssd1 vssd1 vccd1 vccd1 _6729_/A
+ sky130_fd_sc_hd__a32o_1
X_4898_ _4898_/A vssd1 vssd1 vccd1 vccd1 _4900_/B sky130_fd_sc_hd__inv_2
X_7686_ _7711_/A _7711_/B _7685_/X vssd1 vssd1 vccd1 vccd1 _7712_/B sky130_fd_sc_hd__a21o_2
X_6637_ _6637_/A _6663_/B vssd1 vssd1 vccd1 vccd1 _6637_/Y sky130_fd_sc_hd__nand2_1
X_6568_ _8699_/Q _8616_/Q vssd1 vssd1 vccd1 vccd1 _6578_/B sky130_fd_sc_hd__xnor2_4
XFILLER_98_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8307_ _8368_/A _8474_/A vssd1 vssd1 vccd1 vccd1 _8311_/A sky130_fd_sc_hd__or2_1
X_5519_ _5519_/A _5519_/B vssd1 vssd1 vccd1 vccd1 _5525_/A sky130_fd_sc_hd__xnor2_1
X_6499_ _6536_/A _6497_/X _6528_/A _8704_/Q vssd1 vssd1 vccd1 vccd1 _6500_/B sky130_fd_sc_hd__a31o_1
X_8238_ _8238_/A _8238_/B vssd1 vssd1 vccd1 vccd1 _8300_/B sky130_fd_sc_hd__xor2_1
X_8169_ _8378_/A _8242_/B vssd1 vssd1 vccd1 vccd1 _8172_/B sky130_fd_sc_hd__xor2_1
XFILLER_101_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5870_ _5801_/A _5870_/B vssd1 vssd1 vccd1 vccd1 _5870_/X sky130_fd_sc_hd__and2b_1
XFILLER_18_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4821_ _5066_/A _4863_/A _4820_/X vssd1 vssd1 vccd1 vccd1 _5037_/A sky130_fd_sc_hd__o21a_1
X_8752__19 vssd1 vssd1 vccd1 vccd1 _8752__19/HI _8847_/A sky130_fd_sc_hd__conb_1
XFILLER_33_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7540_ _7540_/A _8696_/Q vssd1 vssd1 vccd1 vccd1 _7546_/B sky130_fd_sc_hd__or2_1
X_4752_ _4752_/A _4752_/B vssd1 vssd1 vccd1 vccd1 _4752_/X sky130_fd_sc_hd__or2_1
XFILLER_21_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4683_ _5243_/A vssd1 vssd1 vccd1 vccd1 _5175_/A sky130_fd_sc_hd__clkbuf_2
X_7471_ _7495_/A _7494_/A vssd1 vssd1 vccd1 vccd1 _7505_/A sky130_fd_sc_hd__xnor2_1
X_6422_ _6426_/A _6426_/C vssd1 vssd1 vccd1 vccd1 _6425_/A sky130_fd_sc_hd__and2_1
X_6353_ _6353_/A _6353_/B vssd1 vssd1 vccd1 vccd1 _6354_/B sky130_fd_sc_hd__or2_1
X_5304_ _8635_/Q _8634_/Q _8636_/Q vssd1 vssd1 vccd1 vccd1 _5305_/C sky130_fd_sc_hd__a21o_1
XFILLER_88_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6284_ _6230_/A _6230_/B _6283_/X vssd1 vssd1 vccd1 vccd1 _6289_/A sky130_fd_sc_hd__a21oi_1
XFILLER_88_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5235_ _5202_/D _5226_/X _5234_/X _4960_/A vssd1 vssd1 vccd1 vccd1 _5235_/X sky130_fd_sc_hd__o22a_1
X_8023_ _8023_/A _8023_/B vssd1 vssd1 vccd1 vccd1 _8110_/A sky130_fd_sc_hd__nand2_2
XFILLER_96_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5166_ _5166_/A _5166_/B _5199_/C _5208_/C vssd1 vssd1 vccd1 vccd1 _5166_/X sky130_fd_sc_hd__or4_1
XFILLER_56_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5097_ _5097_/A _5114_/A vssd1 vssd1 vccd1 vccd1 _5109_/B sky130_fd_sc_hd__or2_2
X_8925_ _8925_/A _4445_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[24] sky130_fd_sc_hd__ebufn_8
XFILLER_44_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8856_ _8856_/A _4363_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[25] sky130_fd_sc_hd__ebufn_8
XFILLER_52_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7807_ _8281_/B _7905_/B vssd1 vssd1 vccd1 vccd1 _7903_/C sky130_fd_sc_hd__nor2_1
X_5999_ _5794_/B _6219_/S _5889_/B _5998_/Y vssd1 vssd1 vccd1 vccd1 _6000_/B sky130_fd_sc_hd__a22o_1
XFILLER_12_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7738_ _8620_/Q _8723_/Q vssd1 vssd1 vccd1 vccd1 _7738_/X sky130_fd_sc_hd__or2b_1
X_7669_ _8281_/A _8365_/A vssd1 vssd1 vccd1 vccd1 _7670_/S sky130_fd_sc_hd__or2_1
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5020_ _5035_/A _5194_/C vssd1 vssd1 vccd1 vccd1 _5179_/B sky130_fd_sc_hd__or2_2
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6971_ _7350_/A _7128_/B _7352_/A vssd1 vssd1 vccd1 vccd1 _6973_/B sky130_fd_sc_hd__a21oi_1
X_8710_ _8710_/CLK _8710_/D vssd1 vssd1 vccd1 vccd1 _8710_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5922_ _5922_/A _5922_/B _5922_/C vssd1 vssd1 vccd1 vccd1 _5923_/B sky130_fd_sc_hd__nor3_1
X_8641_ _8681_/CLK _8641_/D vssd1 vssd1 vccd1 vccd1 _8641_/Q sky130_fd_sc_hd__dfxtp_1
X_5853_ _5847_/A _5847_/B _5846_/A vssd1 vssd1 vccd1 vccd1 _5928_/A sky130_fd_sc_hd__o21ai_1
X_8572_ _8572_/A _8576_/B vssd1 vssd1 vccd1 vccd1 _8573_/B sky130_fd_sc_hd__nand2_1
XFILLER_61_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4804_ _4787_/A _4786_/A _4799_/A _4774_/B _4781_/A vssd1 vssd1 vccd1 vccd1 _4804_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_21_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5784_ _5784_/A _6020_/B vssd1 vssd1 vccd1 vccd1 _6204_/B sky130_fd_sc_hd__nand2_2
X_7523_ _7523_/A _7523_/B vssd1 vssd1 vccd1 vccd1 _7523_/X sky130_fd_sc_hd__xor2_1
X_4735_ _4732_/X _4733_/X _4734_/Y vssd1 vssd1 vccd1 vccd1 _8611_/D sky130_fd_sc_hd__o21a_1
XFILLER_21_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7454_ _7454_/A _7454_/B _7454_/C vssd1 vssd1 vccd1 vccd1 _7456_/A sky130_fd_sc_hd__and3_1
X_4666_ _5226_/A vssd1 vssd1 vccd1 vccd1 _5205_/A sky130_fd_sc_hd__clkbuf_2
X_7385_ _7429_/B _7385_/B _7385_/C vssd1 vssd1 vccd1 vccd1 _7387_/A sky130_fd_sc_hd__nor3_1
X_6405_ _8676_/Q _8675_/Q vssd1 vssd1 vccd1 vccd1 _6406_/C sky130_fd_sc_hd__nand2_1
X_4597_ _4597_/A _4597_/B vssd1 vssd1 vccd1 vccd1 _8584_/D sky130_fd_sc_hd__nor2_1
XFILLER_1_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6336_ _6336_/A _6336_/B _6335_/X vssd1 vssd1 vccd1 vccd1 _6336_/X sky130_fd_sc_hd__or3b_1
XFILLER_88_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6267_ _6267_/A _6267_/B vssd1 vssd1 vccd1 vccd1 _6281_/A sky130_fd_sc_hd__xnor2_1
X_5218_ _5218_/A _5218_/B _5218_/C _5218_/D vssd1 vssd1 vccd1 vccd1 _5218_/X sky130_fd_sc_hd__or4_1
XFILLER_69_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6198_ _6198_/A _6198_/B vssd1 vssd1 vccd1 vccd1 _6229_/A sky130_fd_sc_hd__xnor2_4
X_8006_ _8003_/X _8004_/Y _7945_/X _7928_/X vssd1 vssd1 vccd1 vccd1 _8011_/B sky130_fd_sc_hd__a211o_1
X_5149_ _5083_/X _5148_/X _5149_/S vssd1 vssd1 vccd1 vccd1 _5149_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8908_ _8908_/A _4416_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[7] sky130_fd_sc_hd__ebufn_8
X_8839_ _8839_/A _4342_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[8] sky130_fd_sc_hd__ebufn_8
XFILLER_52_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4520_ _5245_/A vssd1 vssd1 vccd1 vccd1 _5199_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_11_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4451_ _4455_/A vssd1 vssd1 vccd1 vccd1 _4451_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7170_ _7170_/A _7170_/B vssd1 vssd1 vccd1 vccd1 _7213_/D sky130_fd_sc_hd__xnor2_1
XFILLER_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4382_ _4382_/A vssd1 vssd1 vccd1 vccd1 _4382_/Y sky130_fd_sc_hd__inv_2
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6121_ _6122_/A _6122_/B vssd1 vssd1 vccd1 vccd1 _6121_/Y sky130_fd_sc_hd__nand2_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6052_ _6048_/A _6052_/B vssd1 vssd1 vccd1 vccd1 _6052_/X sky130_fd_sc_hd__and2b_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5003_ _5016_/A _5227_/D _5208_/C _5245_/D vssd1 vssd1 vccd1 vccd1 _5003_/X sky130_fd_sc_hd__or4_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6954_ _6954_/A _7444_/A vssd1 vssd1 vccd1 vccd1 _6964_/A sky130_fd_sc_hd__and2_1
XFILLER_93_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5905_ _5905_/A _5905_/B vssd1 vssd1 vccd1 vccd1 _5965_/B sky130_fd_sc_hd__xor2_2
X_6885_ _7324_/A _7310_/A vssd1 vssd1 vccd1 vccd1 _7003_/A sky130_fd_sc_hd__nor2_2
X_8624_ _8733_/CLK _8624_/D vssd1 vssd1 vccd1 vccd1 _8624_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5836_ _5943_/A vssd1 vssd1 vccd1 vccd1 _6194_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_22_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5767_ _5767_/A _5767_/B vssd1 vssd1 vccd1 vccd1 _5768_/B sky130_fd_sc_hd__or2_1
X_8555_ _8550_/A _8550_/B _8548_/A vssd1 vssd1 vccd1 vccd1 _8562_/B sky130_fd_sc_hd__a21oi_1
X_4718_ _4718_/A _5080_/B vssd1 vssd1 vccd1 vccd1 _5034_/B sky130_fd_sc_hd__nand2_1
X_7506_ _7509_/B _7505_/Y _7510_/A vssd1 vssd1 vccd1 vccd1 _7506_/X sky130_fd_sc_hd__o21a_1
X_8486_ _8486_/A _8486_/B vssd1 vssd1 vccd1 vccd1 _8492_/A sky130_fd_sc_hd__xnor2_1
X_5698_ _5699_/A _5699_/B vssd1 vssd1 vccd1 vccd1 _5698_/X sky130_fd_sc_hd__or2_1
X_7437_ _7328_/A _7328_/B _7436_/X vssd1 vssd1 vccd1 vccd1 _7441_/A sky130_fd_sc_hd__a21o_1
X_4649_ input2/X vssd1 vssd1 vccd1 vccd1 _5296_/A sky130_fd_sc_hd__clkbuf_2
X_7368_ _7447_/C _7367_/B _7367_/C vssd1 vssd1 vccd1 vccd1 _7373_/B sky130_fd_sc_hd__a21o_1
X_7299_ _7299_/A _7299_/B vssd1 vssd1 vccd1 vccd1 _7391_/A sky130_fd_sc_hd__nor2_1
X_6319_ _6336_/A _6336_/B _6332_/B vssd1 vssd1 vccd1 vccd1 _6319_/X sky130_fd_sc_hd__or3b_1
XFILLER_103_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8788__55 vssd1 vssd1 vccd1 vccd1 _8788__55/HI _8897_/A sky130_fd_sc_hd__conb_1
XFILLER_29_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6670_ _6670_/A _6670_/B vssd1 vssd1 vccd1 vccd1 _7130_/A sky130_fd_sc_hd__nor2_2
XFILLER_50_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5621_ _5621_/A _5621_/B vssd1 vssd1 vccd1 vccd1 _5630_/B sky130_fd_sc_hd__nor2_2
X_8340_ _8415_/A _8341_/B _8413_/B vssd1 vssd1 vccd1 vccd1 _8342_/A sky130_fd_sc_hd__a21oi_1
X_5552_ _5552_/A _5557_/B _5552_/C vssd1 vssd1 vccd1 vccd1 _5556_/A sky130_fd_sc_hd__nand3_1
X_4503_ _8620_/Q vssd1 vssd1 vccd1 vccd1 _7737_/B sky130_fd_sc_hd__buf_2
X_8271_ _8271_/A _8271_/B vssd1 vssd1 vccd1 vccd1 _8271_/Y sky130_fd_sc_hd__nor2_1
X_5483_ _5499_/A _5483_/B vssd1 vssd1 vccd1 vccd1 _5513_/B sky130_fd_sc_hd__xnor2_1
X_4434_ _4437_/A vssd1 vssd1 vccd1 vccd1 _4434_/Y sky130_fd_sc_hd__inv_2
X_7222_ _7188_/Y _7217_/X _7216_/Y _7209_/X vssd1 vssd1 vccd1 vccd1 _7223_/C sky130_fd_sc_hd__o211a_1
XFILLER_104_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4365_ _4369_/A vssd1 vssd1 vccd1 vccd1 _4365_/Y sky130_fd_sc_hd__inv_2
X_7153_ _7157_/A _7157_/B vssd1 vssd1 vccd1 vccd1 _7190_/C sky130_fd_sc_hd__xnor2_1
XFILLER_86_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7084_ _7172_/C _7085_/B _7083_/X vssd1 vssd1 vccd1 vccd1 _7101_/A sky130_fd_sc_hd__a21o_2
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6104_ _6033_/X _6096_/B _6106_/A vssd1 vssd1 vccd1 vccd1 _6113_/A sky130_fd_sc_hd__a21o_1
XFILLER_86_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6035_ _6038_/A _6035_/B vssd1 vssd1 vccd1 vccd1 _6036_/A sky130_fd_sc_hd__xor2_1
XFILLER_100_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7986_ _8066_/A _8071_/A vssd1 vssd1 vccd1 vccd1 _8167_/A sky130_fd_sc_hd__nand2_2
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6937_ _6856_/A _6856_/B _6936_/X vssd1 vssd1 vccd1 vccd1 _6938_/B sky130_fd_sc_hd__o21a_1
XFILLER_25_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6868_ _6868_/A _6779_/B vssd1 vssd1 vccd1 vccd1 _6901_/A sky130_fd_sc_hd__or2b_1
XFILLER_22_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8607_ _8671_/CLK _8607_/D vssd1 vssd1 vccd1 vccd1 _8607_/Q sky130_fd_sc_hd__dfxtp_2
X_5819_ _5819_/A _5819_/B vssd1 vssd1 vccd1 vccd1 _5861_/A sky130_fd_sc_hd__xor2_2
X_6799_ _6724_/A _6798_/Y _6722_/X vssd1 vssd1 vccd1 vccd1 _6801_/A sky130_fd_sc_hd__a21oi_2
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8538_ _7695_/A _7584_/X _8537_/Y vssd1 vssd1 vccd1 vccd1 _8729_/D sky130_fd_sc_hd__o21a_1
X_8469_ _8373_/A _8469_/B vssd1 vssd1 vccd1 vccd1 _8469_/X sky130_fd_sc_hd__and2b_1
XFILLER_89_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7840_ _8515_/C _8205_/A vssd1 vssd1 vccd1 vccd1 _8514_/B sky130_fd_sc_hd__nor2_1
XFILLER_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4983_ _5154_/A _5240_/B _4927_/D _5190_/B vssd1 vssd1 vccd1 vccd1 _4984_/D sky130_fd_sc_hd__a211o_1
XFILLER_63_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7771_ _7771_/A _7771_/B _7771_/C vssd1 vssd1 vccd1 vccd1 _7955_/C sky130_fd_sc_hd__and3_1
X_6722_ _6722_/A _6722_/B _7351_/A vssd1 vssd1 vccd1 vccd1 _6722_/X sky130_fd_sc_hd__and3_1
XFILLER_23_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6653_ _6659_/A _6652_/B _6652_/C vssd1 vssd1 vccd1 vccd1 _6870_/B sky130_fd_sc_hd__a21o_1
X_5604_ _5619_/A _5604_/B vssd1 vssd1 vccd1 vccd1 _5605_/B sky130_fd_sc_hd__nand2_1
X_6584_ _7009_/B vssd1 vssd1 vccd1 vccd1 _7430_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_11_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5535_ _5535_/A _5558_/B _5535_/C vssd1 vssd1 vccd1 vccd1 _5550_/A sky130_fd_sc_hd__and3_1
X_8323_ _8323_/A _8323_/B _8323_/C vssd1 vssd1 vccd1 vccd1 _8324_/B sky130_fd_sc_hd__nor3_1
X_8254_ _8299_/A _8254_/B vssd1 vssd1 vccd1 vccd1 _8256_/C sky130_fd_sc_hd__and2b_1
X_5466_ _5784_/A vssd1 vssd1 vccd1 vccd1 _5892_/A sky130_fd_sc_hd__buf_2
X_7205_ _7213_/B _7128_/B _7275_/A vssd1 vssd1 vccd1 vccd1 _7206_/B sky130_fd_sc_hd__a21oi_1
X_4417_ _4419_/A vssd1 vssd1 vccd1 vccd1 _4417_/Y sky130_fd_sc_hd__inv_2
X_8185_ _8185_/A vssd1 vssd1 vccd1 vccd1 _8499_/A sky130_fd_sc_hd__clkbuf_1
X_5397_ _5397_/A vssd1 vssd1 vccd1 vccd1 _5397_/X sky130_fd_sc_hd__clkbuf_2
X_4348_ _4351_/A vssd1 vssd1 vccd1 vccd1 _4348_/Y sky130_fd_sc_hd__inv_2
X_7136_ _7136_/A _7136_/B vssd1 vssd1 vccd1 vccd1 _7181_/A sky130_fd_sc_hd__xnor2_2
XFILLER_86_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7067_ _7067_/A _7067_/B vssd1 vssd1 vccd1 vccd1 _7211_/A sky130_fd_sc_hd__xor2_2
XFILLER_74_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6018_ _6018_/A _6018_/B vssd1 vssd1 vccd1 vccd1 _6056_/B sky130_fd_sc_hd__xnor2_1
X_8758__25 vssd1 vssd1 vccd1 vccd1 _8758__25/HI _8853_/A sky130_fd_sc_hd__conb_1
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7969_ _8025_/B _7968_/C _7968_/A vssd1 vssd1 vccd1 vccd1 _7976_/B sky130_fd_sc_hd__a21o_1
XFILLER_27_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5320_ _8640_/Q _5322_/C _5308_/X vssd1 vssd1 vccd1 vccd1 _5321_/B sky130_fd_sc_hd__o21ai_1
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5251_ _5096_/A _5206_/X _5216_/X _5221_/X _5250_/X vssd1 vssd1 vccd1 vccd1 _5251_/X
+ sky130_fd_sc_hd__o41a_1
XFILLER_102_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5182_ _5193_/A _5194_/C vssd1 vssd1 vccd1 vccd1 _5183_/C sky130_fd_sc_hd__or2_1
XFILLER_68_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8872_ _8872_/A _4382_/Y vssd1 vssd1 vccd1 vccd1 io_out[9] sky130_fd_sc_hd__ebufn_8
XFILLER_24_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7823_ _7934_/A _7823_/B vssd1 vssd1 vccd1 vccd1 _7825_/B sky130_fd_sc_hd__nand2_1
X_7754_ _8734_/Q _8610_/Q vssd1 vssd1 vccd1 vccd1 _7769_/B sky130_fd_sc_hd__and2b_1
X_4966_ _4966_/A vssd1 vssd1 vccd1 vccd1 _5214_/A sky130_fd_sc_hd__clkbuf_2
X_6705_ _6704_/A _6704_/B _6704_/C vssd1 vssd1 vccd1 vccd1 _7099_/C sky130_fd_sc_hd__a21o_1
X_4897_ _4920_/B _4904_/B vssd1 vssd1 vccd1 vccd1 _5193_/A sky130_fd_sc_hd__nor2_2
XFILLER_22_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7685_ _8730_/Q _8606_/Q vssd1 vssd1 vccd1 vccd1 _7685_/X sky130_fd_sc_hd__and2b_1
X_6636_ _8703_/Q _8620_/Q vssd1 vssd1 vccd1 vccd1 _6663_/B sky130_fd_sc_hd__or2b_1
X_6567_ _7082_/A vssd1 vssd1 vccd1 vccd1 _7128_/A sky130_fd_sc_hd__clkbuf_2
X_8306_ _8367_/A _8306_/B vssd1 vssd1 vccd1 vccd1 _8314_/A sky130_fd_sc_hd__xnor2_2
X_5518_ _5874_/B _5503_/A _5531_/A vssd1 vssd1 vccd1 vccd1 _5521_/C sky130_fd_sc_hd__a21o_1
Xclkbuf_4_1_0_wb_clk_i clkbuf_4_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _8674_/CLK
+ sky130_fd_sc_hd__clkbuf_2
X_6498_ _6498_/A _6536_/B vssd1 vssd1 vccd1 vccd1 _6528_/A sky130_fd_sc_hd__nand2_1
X_8237_ _8237_/A _8237_/B vssd1 vssd1 vccd1 vccd1 _8238_/B sky130_fd_sc_hd__xnor2_2
X_5449_ _8607_/Q _5456_/A vssd1 vssd1 vccd1 vccd1 _5450_/B sky130_fd_sc_hd__and2b_1
XFILLER_87_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8168_ _8515_/B _8166_/X _8069_/B _8167_/Y vssd1 vssd1 vccd1 vccd1 _8242_/B sky130_fd_sc_hd__a31o_1
X_7119_ _7119_/A _7119_/B vssd1 vssd1 vccd1 vccd1 _7120_/B sky130_fd_sc_hd__xnor2_1
XFILLER_59_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8099_ _8265_/A _8265_/B vssd1 vssd1 vccd1 vccd1 _8503_/B sky130_fd_sc_hd__xor2_2
XFILLER_74_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4820_ _4864_/A _4820_/B _4823_/B vssd1 vssd1 vccd1 vccd1 _4820_/X sky130_fd_sc_hd__and3_1
X_4751_ _4660_/A _4660_/B _5087_/A _5634_/B vssd1 vssd1 vccd1 vccd1 _4752_/B sky130_fd_sc_hd__and4bb_1
X_4682_ _5230_/A vssd1 vssd1 vccd1 vccd1 _5243_/A sky130_fd_sc_hd__clkbuf_2
X_7470_ _7493_/A _7493_/B vssd1 vssd1 vccd1 vccd1 _7494_/A sky130_fd_sc_hd__nor2_1
X_6421_ _6421_/A vssd1 vssd1 vccd1 vccd1 _8680_/D sky130_fd_sc_hd__clkbuf_1
X_6352_ _5456_/A _5410_/X _6351_/X _4746_/X vssd1 vssd1 vccd1 vccd1 _8670_/D sky130_fd_sc_hd__o211a_1
X_5303_ _8636_/Q _8635_/Q _8634_/Q vssd1 vssd1 vccd1 vccd1 _5307_/B sky130_fd_sc_hd__and3_1
X_6283_ _6231_/A _6283_/B vssd1 vssd1 vccd1 vccd1 _6283_/X sky130_fd_sc_hd__and2b_1
X_5234_ _5215_/B _5229_/X _5232_/X _5233_/X vssd1 vssd1 vccd1 vccd1 _5234_/X sky130_fd_sc_hd__o22a_1
XFILLER_69_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8022_ _8022_/A _8003_/X vssd1 vssd1 vccd1 vccd1 _8108_/B sky130_fd_sc_hd__or2b_1
X_5165_ _4665_/A _5003_/X _4992_/X _5120_/D _5164_/X vssd1 vssd1 vccd1 vccd1 _5165_/X
+ sky130_fd_sc_hd__o221a_1
X_5096_ _5096_/A _5096_/B _5096_/C _5096_/D vssd1 vssd1 vccd1 vccd1 _5096_/X sky130_fd_sc_hd__or4_1
XFILLER_68_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8924_ _8924_/A _4443_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[23] sky130_fd_sc_hd__ebufn_8
XFILLER_17_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8855_ _8855_/A _4362_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[24] sky130_fd_sc_hd__ebufn_8
XFILLER_71_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7806_ _7836_/A _8065_/B vssd1 vssd1 vccd1 vccd1 _7818_/A sky130_fd_sc_hd__nand2_1
XFILLER_24_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5998_ _5998_/A _6253_/A vssd1 vssd1 vccd1 vccd1 _5998_/Y sky130_fd_sc_hd__nor2_1
X_4949_ _5192_/A _4882_/X vssd1 vssd1 vccd1 vccd1 _5126_/B sky130_fd_sc_hd__or2b_1
XFILLER_33_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7737_ _7618_/A _7737_/B vssd1 vssd1 vccd1 vccd1 _7739_/A sky130_fd_sc_hd__and2b_1
X_7668_ _7798_/B vssd1 vssd1 vccd1 vccd1 _8365_/A sky130_fd_sc_hd__clkbuf_2
X_6619_ _7443_/A _7279_/A vssd1 vssd1 vccd1 vccd1 _6619_/Y sky130_fd_sc_hd__nand2_2
XFILLER_20_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7599_ _7599_/A _7599_/B vssd1 vssd1 vccd1 vccd1 _7599_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_75_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6970_ _7352_/A _7352_/B vssd1 vssd1 vccd1 vccd1 _6973_/A sky130_fd_sc_hd__nor2_1
X_8812__79 vssd1 vssd1 vccd1 vccd1 _8812__79/HI _8921_/A sky130_fd_sc_hd__conb_1
XFILLER_93_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5921_ _5922_/A _5922_/B _5922_/C vssd1 vssd1 vccd1 vccd1 _5923_/A sky130_fd_sc_hd__o21a_1
XFILLER_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8640_ _8681_/CLK _8640_/D vssd1 vssd1 vccd1 vccd1 _8640_/Q sky130_fd_sc_hd__dfxtp_1
X_5852_ _6058_/A _6058_/B vssd1 vssd1 vccd1 vccd1 _6060_/B sky130_fd_sc_hd__nor2_1
X_4803_ _4801_/B _4720_/A _4715_/B _4732_/X _4802_/Y vssd1 vssd1 vccd1 vccd1 _4803_/X
+ sky130_fd_sc_hd__a41o_1
X_8571_ _8571_/A _8571_/B vssd1 vssd1 vccd1 vccd1 _8576_/B sky130_fd_sc_hd__or2_1
X_5783_ _5708_/A _5795_/A _5777_/B _5574_/A vssd1 vssd1 vccd1 vccd1 _5798_/A sky130_fd_sc_hd__a22o_1
X_7522_ _7514_/A _7526_/B _7515_/Y vssd1 vssd1 vccd1 vccd1 _7523_/B sky130_fd_sc_hd__a21o_1
X_4734_ _4730_/B _4732_/X _4727_/A vssd1 vssd1 vccd1 vccd1 _4734_/Y sky130_fd_sc_hd__a21boi_1
X_7453_ _7378_/C _7378_/Y _7451_/Y _7452_/Y vssd1 vssd1 vccd1 vccd1 _7457_/A sky130_fd_sc_hd__o31ai_1
X_4665_ _4665_/A vssd1 vssd1 vccd1 vccd1 _5028_/B sky130_fd_sc_hd__clkbuf_2
X_7384_ _7018_/B _7018_/C _7018_/A vssd1 vssd1 vccd1 vccd1 _7385_/C sky130_fd_sc_hd__o21ba_1
X_6404_ _6457_/B vssd1 vssd1 vccd1 vccd1 _6406_/B sky130_fd_sc_hd__clkbuf_2
X_4596_ _8584_/Q _4598_/C _4595_/X vssd1 vssd1 vccd1 vccd1 _4597_/B sky130_fd_sc_hd__o21ai_1
X_6335_ _6295_/A _6296_/X _6335_/S vssd1 vssd1 vccd1 vccd1 _6335_/X sky130_fd_sc_hd__mux2_1
XFILLER_103_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6266_ _6266_/A _6266_/B vssd1 vssd1 vccd1 vccd1 _6267_/B sky130_fd_sc_hd__xnor2_1
X_8005_ _7945_/X _7928_/X _8003_/X _8004_/Y vssd1 vssd1 vccd1 vccd1 _8021_/A sky130_fd_sc_hd__o211ai_2
X_5217_ _5173_/A _5169_/A _5109_/C _5173_/Y _5196_/B vssd1 vssd1 vccd1 vccd1 _5218_/C
+ sky130_fd_sc_hd__o32a_1
XFILLER_57_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6197_ _6197_/A _6262_/A vssd1 vssd1 vccd1 vccd1 _6198_/B sky130_fd_sc_hd__xnor2_2
XFILLER_96_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5148_ _5080_/Y _5096_/X _5125_/X _5147_/X vssd1 vssd1 vccd1 vccd1 _5148_/X sky130_fd_sc_hd__a31o_1
X_5079_ _5079_/A _5248_/A vssd1 vssd1 vccd1 vccd1 _5080_/A sky130_fd_sc_hd__nor2_1
XFILLER_17_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8907_ _8907_/A _4413_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[6] sky130_fd_sc_hd__ebufn_8
XFILLER_71_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8838_ _8838_/A _4341_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[7] sky130_fd_sc_hd__ebufn_8
XFILLER_12_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4450_ _4456_/A vssd1 vssd1 vccd1 vccd1 _4455_/A sky130_fd_sc_hd__buf_2
XFILLER_7_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4381_ _4382_/A vssd1 vssd1 vccd1 vccd1 _4381_/Y sky130_fd_sc_hd__inv_2
X_6120_ _6120_/A _6120_/B vssd1 vssd1 vccd1 vccd1 _6133_/A sky130_fd_sc_hd__or2_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6051_ _6051_/A _6055_/B vssd1 vssd1 vccd1 vccd1 _6085_/B sky130_fd_sc_hd__xnor2_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5002_ _5186_/A _5002_/B vssd1 vssd1 vccd1 vccd1 _5208_/C sky130_fd_sc_hd__or2_2
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6953_ _7327_/A vssd1 vssd1 vccd1 vccd1 _7444_/A sky130_fd_sc_hd__clkbuf_2
X_6884_ _6884_/A _7004_/A vssd1 vssd1 vccd1 vccd1 _6951_/A sky130_fd_sc_hd__or2b_1
X_5904_ _5904_/A _5904_/B vssd1 vssd1 vccd1 vccd1 _5905_/B sky130_fd_sc_hd__xor2_2
XFILLER_22_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8623_ _8733_/CLK _8623_/D vssd1 vssd1 vccd1 vccd1 _8623_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5835_ _6182_/A _5909_/B vssd1 vssd1 vccd1 vccd1 _5838_/B sky130_fd_sc_hd__xor2_1
X_8554_ _8563_/A _8554_/B vssd1 vssd1 vccd1 vccd1 _8556_/A sky130_fd_sc_hd__or2_1
X_5766_ _5767_/A _5767_/B vssd1 vssd1 vccd1 vccd1 _5847_/A sky130_fd_sc_hd__nand2_1
X_4717_ _4714_/A _4716_/A _4716_/Y _4672_/X vssd1 vssd1 vccd1 vccd1 _8607_/D sky130_fd_sc_hd__o211a_1
X_7505_ _7505_/A _7505_/B vssd1 vssd1 vccd1 vccd1 _7505_/Y sky130_fd_sc_hd__nor2_1
X_8485_ _8485_/A _8485_/B vssd1 vssd1 vccd1 vccd1 _8486_/B sky130_fd_sc_hd__xnor2_1
X_5697_ _5584_/A _5584_/B _5696_/X vssd1 vssd1 vccd1 vccd1 _5727_/A sky130_fd_sc_hd__a21oi_2
X_7436_ _7444_/A _7436_/B vssd1 vssd1 vccd1 vccd1 _7436_/X sky130_fd_sc_hd__and2_1
X_4648_ _8601_/Q _4648_/B vssd1 vssd1 vccd1 vccd1 _4648_/Y sky130_fd_sc_hd__nand2_1
XFILLER_30_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7367_ _7447_/C _7367_/B _7367_/C vssd1 vssd1 vccd1 vccd1 _7447_/D sky130_fd_sc_hd__nand3_1
X_4579_ _4647_/A _8601_/Q vssd1 vssd1 vccd1 vccd1 _5434_/B sky130_fd_sc_hd__or2b_1
XFILLER_1_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7298_ _7475_/A _7479_/B _7475_/C _7484_/B _7297_/X vssd1 vssd1 vccd1 vccd1 _7489_/S
+ sky130_fd_sc_hd__a41o_1
XFILLER_1_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6318_ _6134_/A _5831_/X _6316_/Y _6317_/Y _6321_/A vssd1 vssd1 vccd1 vccd1 _6332_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6249_ _6249_/A _6249_/B vssd1 vssd1 vccd1 vccd1 _6250_/B sky130_fd_sc_hd__xnor2_2
XFILLER_49_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_4_14_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8715_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5620_ _7737_/B _8662_/Q vssd1 vssd1 vccd1 vccd1 _5621_/A sky130_fd_sc_hd__and2b_1
X_5551_ _5550_/A _5550_/B _5549_/Y vssd1 vssd1 vccd1 vccd1 _5552_/C sky130_fd_sc_hd__o21bai_1
X_4502_ _4765_/A _4790_/A vssd1 vssd1 vccd1 vccd1 _4786_/B sky130_fd_sc_hd__and2_1
XFILLER_8_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8270_ _8499_/A _8501_/B _8499_/B vssd1 vssd1 vccd1 vccd1 _8496_/C sky130_fd_sc_hd__o21ai_1
X_7221_ _7215_/A _7219_/Y _7220_/Y vssd1 vssd1 vccd1 vccd1 _7223_/B sky130_fd_sc_hd__o21a_1
X_5482_ _5566_/A _5784_/A _5479_/Y _6020_/B vssd1 vssd1 vccd1 vccd1 _5483_/B sky130_fd_sc_hd__o211a_1
X_4433_ _4437_/A vssd1 vssd1 vccd1 vccd1 _4433_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4364_ _4370_/A vssd1 vssd1 vccd1 vccd1 _4369_/A sky130_fd_sc_hd__clkbuf_2
X_7152_ _7152_/A _7152_/B vssd1 vssd1 vccd1 vccd1 _7157_/B sky130_fd_sc_hd__xnor2_1
XFILLER_98_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7083_ _7169_/A _7083_/B _7170_/A vssd1 vssd1 vccd1 vccd1 _7083_/X sky130_fd_sc_hd__and3_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6103_ _5831_/X _6095_/A _6101_/A _6102_/X _6097_/B vssd1 vssd1 vccd1 vccd1 _6106_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_100_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6034_ _6096_/A _6034_/B _6033_/X vssd1 vssd1 vccd1 vccd1 _6036_/B sky130_fd_sc_hd__or3b_2
XFILLER_100_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7985_ _7919_/A _7985_/B vssd1 vssd1 vccd1 vccd1 _7993_/B sky130_fd_sc_hd__and2b_1
X_6936_ _6856_/A _6856_/B _6831_/Y vssd1 vssd1 vccd1 vccd1 _6936_/X sky130_fd_sc_hd__a21bo_1
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6867_ _6819_/A _6819_/B _6790_/A vssd1 vssd1 vccd1 vccd1 _6948_/A sky130_fd_sc_hd__a21o_1
X_6798_ _6876_/B _6972_/C _7074_/C _6774_/S vssd1 vssd1 vccd1 vccd1 _6798_/Y sky130_fd_sc_hd__o31ai_2
X_8606_ _8714_/CLK _8606_/D vssd1 vssd1 vccd1 vccd1 _8606_/Q sky130_fd_sc_hd__dfxtp_4
X_5818_ _5943_/A _5970_/A _6193_/B _5817_/Y vssd1 vssd1 vccd1 vccd1 _5819_/B sky130_fd_sc_hd__o31a_1
XFILLER_10_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5749_ _5838_/A _5748_/X vssd1 vssd1 vccd1 vccd1 _5751_/B sky130_fd_sc_hd__or2b_1
XFILLER_10_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8537_ _7695_/A _8574_/A _4785_/A vssd1 vssd1 vccd1 vccd1 _8537_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_41_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8468_ _8377_/A _8377_/B _8378_/B _8378_/A vssd1 vssd1 vccd1 vccd1 _8479_/A sky130_fd_sc_hd__a2bb2o_1
X_8739__6 vssd1 vssd1 vccd1 vccd1 _8739__6/HI _8834_/A sky130_fd_sc_hd__conb_1
X_7419_ _7340_/A _7419_/B vssd1 vssd1 vccd1 vccd1 _7419_/X sky130_fd_sc_hd__and2b_1
X_8399_ _8399_/A _8399_/B vssd1 vssd1 vccd1 vccd1 _8400_/B sky130_fd_sc_hd__xnor2_1
XFILLER_104_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4982_ _5185_/B _5175_/B _5155_/A vssd1 vssd1 vccd1 vccd1 _4984_/C sky130_fd_sc_hd__o21a_1
XFILLER_23_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7770_ _7759_/A _7759_/B _7769_/X vssd1 vssd1 vccd1 vccd1 _7771_/C sky130_fd_sc_hd__a21o_1
X_6721_ _6688_/X _6689_/X _6657_/A vssd1 vssd1 vccd1 vccd1 _7351_/A sky130_fd_sc_hd__a21o_1
X_6652_ _6659_/A _6652_/B _6652_/C vssd1 vssd1 vccd1 vccd1 _6870_/A sky130_fd_sc_hd__nand3_1
X_5603_ _5603_/A vssd1 vssd1 vccd1 vccd1 _5604_/B sky130_fd_sc_hd__inv_2
X_6583_ _6614_/A vssd1 vssd1 vccd1 vccd1 _7009_/B sky130_fd_sc_hd__clkbuf_2
X_8322_ _8323_/B _8323_/C _8323_/A vssd1 vssd1 vccd1 vccd1 _8324_/A sky130_fd_sc_hd__o21a_1
XFILLER_11_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5534_ _5533_/A _5533_/B _5532_/X vssd1 vssd1 vccd1 vccd1 _5535_/C sky130_fd_sc_hd__o21bai_1
X_8253_ _8253_/A _8253_/B vssd1 vssd1 vccd1 vccd1 _8254_/B sky130_fd_sc_hd__nand2_1
X_5465_ _5874_/B _5705_/A vssd1 vssd1 vccd1 vccd1 _5784_/A sky130_fd_sc_hd__nand2_2
X_7204_ _7172_/B _7172_/C _7454_/A vssd1 vssd1 vccd1 vccd1 _7234_/B sky130_fd_sc_hd__o21ai_1
X_4416_ _4419_/A vssd1 vssd1 vccd1 vccd1 _4416_/Y sky130_fd_sc_hd__inv_2
X_8184_ _8266_/A _8266_/B vssd1 vssd1 vccd1 vccd1 _8185_/A sky130_fd_sc_hd__and2_1
X_7135_ _7135_/A _7135_/B vssd1 vssd1 vccd1 vccd1 _7136_/A sky130_fd_sc_hd__xnor2_1
X_5396_ _5396_/A vssd1 vssd1 vccd1 vccd1 _8657_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4347_ _4351_/A vssd1 vssd1 vccd1 vccd1 _4347_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7066_ _7065_/X _6836_/A _7059_/Y vssd1 vssd1 vccd1 vccd1 _7067_/B sky130_fd_sc_hd__o21ba_1
XFILLER_59_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6017_ _6312_/A _6236_/B vssd1 vssd1 vccd1 vccd1 _6302_/A sky130_fd_sc_hd__and2_1
XFILLER_27_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7968_ _7968_/A _8025_/B _7968_/C vssd1 vssd1 vccd1 vccd1 _8024_/A sky130_fd_sc_hd__nand3_1
XFILLER_42_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6919_ _6919_/A _7025_/B vssd1 vssd1 vccd1 vccd1 _6920_/B sky130_fd_sc_hd__xnor2_1
XFILLER_52_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7899_ _7945_/A _7945_/B _7945_/C vssd1 vssd1 vccd1 vccd1 _7928_/A sky130_fd_sc_hd__nand3_1
XFILLER_10_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5250_ _5064_/A _5235_/X _5249_/X _4710_/A vssd1 vssd1 vccd1 vccd1 _5250_/X sky130_fd_sc_hd__a211o_1
XFILLER_5_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5181_ _5186_/A _5227_/B _5179_/X _5180_/X vssd1 vssd1 vccd1 vccd1 _5181_/X sky130_fd_sc_hd__o31a_1
XFILLER_68_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8871_ _8871_/A _4381_/Y vssd1 vssd1 vccd1 vccd1 io_out[8] sky130_fd_sc_hd__ebufn_8
XFILLER_83_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7822_ _7822_/A _7822_/B vssd1 vssd1 vccd1 vccd1 _7823_/B sky130_fd_sc_hd__nand2_1
X_4965_ _5131_/A _4965_/B vssd1 vssd1 vccd1 vccd1 _5172_/A sky130_fd_sc_hd__or2_1
X_7753_ _8610_/Q _8734_/Q vssd1 vssd1 vccd1 vccd1 _7775_/A sky130_fd_sc_hd__and2b_1
X_6704_ _6704_/A _6704_/B _6704_/C vssd1 vssd1 vccd1 vccd1 _7099_/B sky130_fd_sc_hd__nand3_4
X_4896_ _4896_/A _5047_/B vssd1 vssd1 vccd1 vccd1 _5169_/A sky130_fd_sc_hd__nor2_2
X_7684_ _8730_/Q _8606_/Q vssd1 vssd1 vccd1 vccd1 _7711_/B sky130_fd_sc_hd__xnor2_4
X_6635_ _6637_/A _6635_/B vssd1 vssd1 vccd1 vccd1 _6652_/C sky130_fd_sc_hd__and2_1
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6566_ _6588_/A _6588_/B vssd1 vssd1 vccd1 vccd1 _7082_/A sky130_fd_sc_hd__and2_1
X_8305_ _8304_/A _8368_/B _8304_/Y _8071_/A vssd1 vssd1 vccd1 vccd1 _8306_/B sky130_fd_sc_hd__o22a_1
X_5517_ _5517_/A _5998_/A vssd1 vssd1 vccd1 vccd1 _5531_/A sky130_fd_sc_hd__nor2_2
X_6497_ _6509_/A _8698_/Q _6526_/B _6515_/A _6521_/A vssd1 vssd1 vccd1 vccd1 _6497_/X
+ sky130_fd_sc_hd__a2111o_1
X_8236_ _8345_/B _8236_/B vssd1 vssd1 vccd1 vccd1 _8237_/B sky130_fd_sc_hd__nand2_1
X_5448_ _8670_/Q _8607_/Q vssd1 vssd1 vccd1 vccd1 _5450_/A sky130_fd_sc_hd__and2b_1
X_8818__85 vssd1 vssd1 vccd1 vccd1 _8818__85/HI _8927_/A sky130_fd_sc_hd__conb_1
X_8167_ _8167_/A _8291_/A vssd1 vssd1 vccd1 vccd1 _8167_/Y sky130_fd_sc_hd__nor2_1
X_5379_ _5426_/B vssd1 vssd1 vccd1 vccd1 _5425_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_101_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7118_ _7162_/A _7162_/B _7117_/X vssd1 vssd1 vccd1 vccd1 _7120_/A sky130_fd_sc_hd__a21o_1
X_8098_ _8098_/A _8098_/B vssd1 vssd1 vccd1 vccd1 _8265_/B sky130_fd_sc_hd__xor2_2
X_7049_ _7046_/X _7047_/X _7299_/A _7045_/Y vssd1 vssd1 vccd1 vccd1 _7299_/B sky130_fd_sc_hd__a211oi_2
XFILLER_74_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4750_ _4848_/A _4848_/B _4834_/C _4839_/A vssd1 vssd1 vccd1 vccd1 _5087_/A sky130_fd_sc_hd__and4b_2
XFILLER_14_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4681_ _5185_/A vssd1 vssd1 vccd1 vccd1 _5230_/A sky130_fd_sc_hd__clkbuf_2
X_6420_ _6426_/C _6420_/B _6457_/B vssd1 vssd1 vccd1 vccd1 _6421_/A sky130_fd_sc_hd__and3b_1
X_6351_ _6355_/B _6350_/Y _4581_/B vssd1 vssd1 vccd1 vccd1 _6351_/X sky130_fd_sc_hd__a21o_1
X_5302_ _5302_/A vssd1 vssd1 vccd1 vccd1 _8635_/D sky130_fd_sc_hd__clkbuf_1
X_6282_ _6282_/A _6282_/B vssd1 vssd1 vccd1 vccd1 _6290_/A sky130_fd_sc_hd__xnor2_4
X_5233_ _8604_/Q _5233_/B _5233_/C vssd1 vssd1 vccd1 vccd1 _5233_/X sky130_fd_sc_hd__or3_1
X_8021_ _8021_/A _8021_/B vssd1 vssd1 vccd1 vccd1 _8106_/B sky130_fd_sc_hd__nand2_1
XFILLER_102_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5164_ _5192_/B _5238_/C _5164_/C _5164_/D vssd1 vssd1 vccd1 vccd1 _5164_/X sky130_fd_sc_hd__or4_1
XFILLER_68_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5095_ _5053_/A _5245_/B _5090_/X _5091_/X _5094_/X vssd1 vssd1 vccd1 vccd1 _5096_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_83_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8923_ _8923_/A _4442_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[22] sky130_fd_sc_hd__ebufn_8
XFILLER_71_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8854_ _8854_/A _4361_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[23] sky130_fd_sc_hd__ebufn_8
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7805_ _7805_/A vssd1 vssd1 vccd1 vccd1 _8065_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_24_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5997_ _5997_/A vssd1 vssd1 vccd1 vccd1 _6253_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_33_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4948_ _4990_/A _4948_/B vssd1 vssd1 vccd1 vccd1 _5240_/B sky130_fd_sc_hd__nor2_2
X_7736_ _7736_/A _8515_/B _7833_/B vssd1 vssd1 vccd1 vccd1 _7831_/C sky130_fd_sc_hd__and3_1
X_4879_ _4879_/A _4879_/B vssd1 vssd1 vccd1 vccd1 _5115_/A sky130_fd_sc_hd__nor2_2
X_7667_ _7988_/A vssd1 vssd1 vccd1 vccd1 _7798_/B sky130_fd_sc_hd__clkbuf_2
X_6618_ _6835_/A _7009_/B vssd1 vssd1 vccd1 vccd1 _7279_/A sky130_fd_sc_hd__nor2_2
XFILLER_20_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7598_ _7630_/A _7592_/B _7591_/A vssd1 vssd1 vccd1 vccd1 _7599_/B sky130_fd_sc_hd__o21a_1
X_6549_ _7516_/A _7695_/B vssd1 vssd1 vccd1 vccd1 _6593_/B sky130_fd_sc_hd__nand2_1
X_8219_ _7728_/A _8331_/A _8220_/B _8120_/B _8203_/B vssd1 vssd1 vccd1 vccd1 _8319_/A
+ sky130_fd_sc_hd__a32o_1
XFILLER_58_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5920_ _5964_/A _5920_/B vssd1 vssd1 vccd1 vccd1 _5922_/C sky130_fd_sc_hd__and2b_1
XFILLER_46_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5851_ _5851_/A _5851_/B vssd1 vssd1 vccd1 vccd1 _6058_/B sky130_fd_sc_hd__xnor2_1
X_4802_ _4802_/A vssd1 vssd1 vccd1 vccd1 _4802_/Y sky130_fd_sc_hd__inv_2
X_8570_ _8571_/A _8571_/B vssd1 vssd1 vccd1 vccd1 _8572_/A sky130_fd_sc_hd__nand2_1
X_5782_ _5992_/A _5782_/B vssd1 vssd1 vccd1 vccd1 _5790_/A sky130_fd_sc_hd__xnor2_1
XFILLER_34_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7521_ _7521_/A _7521_/B vssd1 vssd1 vccd1 vccd1 _7523_/A sky130_fd_sc_hd__nor2_1
X_4733_ _4478_/X _4730_/B _4733_/S vssd1 vssd1 vccd1 vccd1 _4733_/X sky130_fd_sc_hd__mux2_1
X_7452_ _7378_/C _7378_/Y _7451_/Y vssd1 vssd1 vccd1 vccd1 _7452_/Y sky130_fd_sc_hd__o21ai_1
X_6403_ input2/X _6403_/B vssd1 vssd1 vccd1 vccd1 _6457_/B sky130_fd_sc_hd__and2_1
X_4664_ _5226_/B _4923_/A vssd1 vssd1 vccd1 vccd1 _4665_/A sky130_fd_sc_hd__nand2_2
X_7383_ _7429_/A _7382_/C _7382_/A vssd1 vssd1 vccd1 vccd1 _7385_/B sky130_fd_sc_hd__o21a_1
X_4595_ _4645_/B vssd1 vssd1 vccd1 vccd1 _4595_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6334_ _6324_/X _6333_/X _6325_/X _8666_/Q vssd1 vssd1 vccd1 vccd1 _8666_/D sky130_fd_sc_hd__o2bb2a_1
XFILLER_103_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6265_ _6265_/A _6265_/B vssd1 vssd1 vccd1 vccd1 _6266_/B sky130_fd_sc_hd__xnor2_1
XFILLER_103_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5216_ _4916_/A _5196_/B _5211_/X _5215_/X _5080_/B vssd1 vssd1 vccd1 vccd1 _5216_/X
+ sky130_fd_sc_hd__o311a_1
X_8004_ _8022_/A _8003_/B _8003_/C vssd1 vssd1 vccd1 vccd1 _8004_/Y sky130_fd_sc_hd__o21ai_1
X_6196_ _6196_/A _6255_/B vssd1 vssd1 vccd1 vccd1 _6262_/A sky130_fd_sc_hd__xnor2_2
X_5147_ _5096_/B _5146_/X _5056_/A vssd1 vssd1 vccd1 vccd1 _5147_/X sky130_fd_sc_hd__o21a_1
XFILLER_69_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5078_ _5248_/A _5193_/A _5078_/C _5078_/D vssd1 vssd1 vccd1 vccd1 _5078_/X sky130_fd_sc_hd__or4_1
XFILLER_84_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8906_ _8906_/A _4415_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[5] sky130_fd_sc_hd__ebufn_8
XFILLER_44_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8837_ _8837_/A _4340_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[6] sky130_fd_sc_hd__ebufn_8
XFILLER_44_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7719_ _7750_/A _7750_/B vssd1 vssd1 vccd1 vccd1 _7734_/A sky130_fd_sc_hd__xnor2_1
XFILLER_100_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8699_ _8733_/CLK _8699_/D vssd1 vssd1 vccd1 vccd1 _8699_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4380_ _4382_/A vssd1 vssd1 vccd1 vccd1 _4380_/Y sky130_fd_sc_hd__clkinv_4
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6050_ _5767_/A _6049_/Y _5687_/A _5687_/B vssd1 vssd1 vccd1 vccd1 _6055_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5001_ _5037_/A vssd1 vssd1 vccd1 vccd1 _5186_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6952_ _6952_/A _6952_/B vssd1 vssd1 vccd1 vccd1 _6952_/Y sky130_fd_sc_hd__nand2_1
XFILLER_81_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6883_ _6883_/A _6883_/B vssd1 vssd1 vccd1 vccd1 _6952_/A sky130_fd_sc_hd__xor2_2
X_5903_ _5903_/A _5903_/B vssd1 vssd1 vccd1 vccd1 _5904_/B sky130_fd_sc_hd__xnor2_2
X_8622_ _8734_/CLK _8622_/D vssd1 vssd1 vccd1 vccd1 _8622_/Q sky130_fd_sc_hd__dfxtp_1
X_5834_ _5831_/X _5953_/A _5745_/B _5833_/Y vssd1 vssd1 vccd1 vccd1 _5909_/B sky130_fd_sc_hd__a31o_1
X_8553_ _8553_/A _8571_/B vssd1 vssd1 vccd1 vccd1 _8554_/B sky130_fd_sc_hd__nor2_1
X_5765_ _5924_/A _5765_/B vssd1 vssd1 vccd1 vccd1 _5767_/B sky130_fd_sc_hd__nor2_1
X_4716_ _4716_/A _5149_/S vssd1 vssd1 vccd1 vccd1 _4716_/Y sky130_fd_sc_hd__nand2_1
X_7504_ _7505_/A _7505_/B vssd1 vssd1 vccd1 vccd1 _7509_/B sky130_fd_sc_hd__and2_1
X_8484_ _8484_/A _8484_/B vssd1 vssd1 vccd1 vccd1 _8485_/B sky130_fd_sc_hd__xnor2_1
X_5696_ _5583_/A _5696_/B vssd1 vssd1 vccd1 vccd1 _5696_/X sky130_fd_sc_hd__and2b_1
X_7435_ _7280_/A _7434_/B _7454_/C _7434_/X vssd1 vssd1 vccd1 vccd1 _7459_/A sky130_fd_sc_hd__o31a_1
X_4647_ _4647_/A vssd1 vssd1 vccd1 vccd1 _5389_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7366_ _7366_/A _7366_/B vssd1 vssd1 vccd1 vccd1 _7367_/C sky130_fd_sc_hd__nand2_1
XFILLER_89_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6317_ _6134_/A _6134_/B _5941_/X vssd1 vssd1 vccd1 vccd1 _6317_/Y sky130_fd_sc_hd__o21bai_1
X_4578_ _4587_/A _4578_/B _4578_/C vssd1 vssd1 vccd1 vccd1 _4647_/A sky130_fd_sc_hd__nor3_1
XFILLER_103_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7297_ _7296_/A _7202_/A _7296_/B vssd1 vssd1 vccd1 vccd1 _7297_/X sky130_fd_sc_hd__o21ba_1
X_6248_ _5981_/B _6246_/Y _6247_/Y vssd1 vssd1 vccd1 vccd1 _6249_/B sky130_fd_sc_hd__o21a_1
X_6179_ _5957_/A _6179_/B vssd1 vssd1 vccd1 vccd1 _6179_/X sky130_fd_sc_hd__and2b_1
XFILLER_57_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8779__46 vssd1 vssd1 vccd1 vccd1 _8779__46/HI _8888_/A sky130_fd_sc_hd__conb_1
XFILLER_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5550_ _5550_/A _5550_/B _5549_/Y vssd1 vssd1 vccd1 vccd1 _5557_/B sky130_fd_sc_hd__or3b_1
X_4501_ _4781_/A _4799_/A _4808_/A vssd1 vssd1 vccd1 vccd1 _4790_/A sky130_fd_sc_hd__and3_2
XFILLER_8_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5481_ _5873_/A _5481_/B vssd1 vssd1 vccd1 vccd1 _6020_/B sky130_fd_sc_hd__nand2_2
X_7220_ _7220_/A _7220_/B vssd1 vssd1 vccd1 vccd1 _7220_/Y sky130_fd_sc_hd__nand2_1
X_4432_ _4432_/A vssd1 vssd1 vccd1 vccd1 _4437_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_104_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4363_ _4363_/A vssd1 vssd1 vccd1 vccd1 _4363_/Y sky130_fd_sc_hd__inv_2
X_7151_ _7151_/A _7151_/B vssd1 vssd1 vccd1 vccd1 _7152_/B sky130_fd_sc_hd__xnor2_1
XFILLER_6_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7082_ _7082_/A _7350_/B vssd1 vssd1 vccd1 vccd1 _7170_/A sky130_fd_sc_hd__nor2_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6102_ _6122_/A _6122_/B vssd1 vssd1 vccd1 vccd1 _6102_/X sky130_fd_sc_hd__and2_1
XFILLER_98_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6033_ _6033_/A _6033_/B vssd1 vssd1 vccd1 vccd1 _6033_/X sky130_fd_sc_hd__and2_1
XFILLER_39_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7984_ _7914_/A _7984_/B vssd1 vssd1 vccd1 vccd1 _8078_/A sky130_fd_sc_hd__and2b_1
X_6935_ _6935_/A _6935_/B vssd1 vssd1 vccd1 vccd1 _7023_/B sky130_fd_sc_hd__xor2_1
XFILLER_81_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8793__60 vssd1 vssd1 vccd1 vccd1 _8793__60/HI _8902_/A sky130_fd_sc_hd__conb_1
XFILLER_41_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6866_ _7115_/A _7115_/B _6865_/X vssd1 vssd1 vccd1 vccd1 _6944_/A sky130_fd_sc_hd__a21o_1
XFILLER_34_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6797_ _6797_/A _7102_/B vssd1 vssd1 vccd1 vccd1 _6802_/A sky130_fd_sc_hd__nor2_1
X_8605_ _8714_/CLK _8605_/D vssd1 vssd1 vccd1 vccd1 _8605_/Q sky130_fd_sc_hd__dfxtp_4
X_5817_ _5943_/A _5970_/A _5816_/B vssd1 vssd1 vccd1 vccd1 _5817_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_10_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5748_ _5945_/A _5747_/B _5747_/D _5747_/C vssd1 vssd1 vccd1 vccd1 _5748_/X sky130_fd_sc_hd__a31o_1
X_8536_ _4771_/X _8520_/X _8534_/X _8535_/Y vssd1 vssd1 vccd1 vccd1 _8728_/D sky130_fd_sc_hd__a31oi_1
XFILLER_41_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5679_ _5680_/A _5680_/B vssd1 vssd1 vccd1 vccd1 _5692_/B sky130_fd_sc_hd__nand2_1
X_8467_ _8467_/A _8467_/B vssd1 vssd1 vccd1 vccd1 _8485_/A sky130_fd_sc_hd__xnor2_1
X_7418_ _7418_/A _7418_/B vssd1 vssd1 vccd1 vccd1 _7423_/A sky130_fd_sc_hd__xnor2_1
X_8398_ _8124_/A _7716_/X _8450_/A vssd1 vssd1 vccd1 vccd1 _8401_/A sky130_fd_sc_hd__a21oi_1
X_7349_ _7349_/A vssd1 vssd1 vccd1 vccd1 _7454_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4981_ _5214_/A _5245_/B _5238_/B vssd1 vssd1 vccd1 vccd1 _5175_/C sky130_fd_sc_hd__or3_2
X_6720_ _6625_/X _6688_/X _6689_/X _6876_/A _7075_/A vssd1 vssd1 vccd1 vccd1 _6722_/A
+ sky130_fd_sc_hd__a311oi_1
XFILLER_16_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6651_ _7103_/A _6651_/B vssd1 vssd1 vccd1 vccd1 _7099_/A sky130_fd_sc_hd__xor2_1
X_6582_ _6593_/A _6582_/B vssd1 vssd1 vccd1 vccd1 _6614_/A sky130_fd_sc_hd__xnor2_2
X_5602_ _8661_/Q _7652_/B vssd1 vssd1 vccd1 vccd1 _5603_/A sky130_fd_sc_hd__and2b_1
X_5533_ _5533_/A _5533_/B _5532_/X vssd1 vssd1 vccd1 vccd1 _5558_/B sky130_fd_sc_hd__or3b_1
X_8321_ _8321_/A _8321_/B vssd1 vssd1 vccd1 vccd1 _8323_/B sky130_fd_sc_hd__nor2_1
X_8252_ _8253_/A _8253_/B vssd1 vssd1 vccd1 vccd1 _8299_/A sky130_fd_sc_hd__nor2_1
X_5464_ _5477_/A _5477_/B vssd1 vssd1 vccd1 vccd1 _5705_/A sky130_fd_sc_hd__xor2_1
X_7203_ _7203_/A _7203_/B vssd1 vssd1 vccd1 vccd1 _7230_/A sky130_fd_sc_hd__xor2_1
X_8183_ _8186_/A _8183_/B vssd1 vssd1 vccd1 vccd1 _8266_/B sky130_fd_sc_hd__xnor2_1
X_5395_ _5397_/A _5398_/A _5615_/A vssd1 vssd1 vccd1 vccd1 _5396_/A sky130_fd_sc_hd__mux2_1
X_4415_ _4419_/A vssd1 vssd1 vccd1 vccd1 _4415_/Y sky130_fd_sc_hd__inv_2
X_4346_ _4370_/A vssd1 vssd1 vccd1 vccd1 _4351_/A sky130_fd_sc_hd__clkbuf_2
X_7134_ _7173_/A _7173_/B _7133_/X vssd1 vssd1 vccd1 vccd1 _7141_/A sky130_fd_sc_hd__a21o_1
XFILLER_101_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7065_ _7065_/A _7430_/B vssd1 vssd1 vccd1 vccd1 _7065_/X sky130_fd_sc_hd__or2_1
X_6016_ _6061_/A _6016_/B vssd1 vssd1 vccd1 vccd1 _6236_/B sky130_fd_sc_hd__nand2_1
XFILLER_27_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7967_ _8025_/A _7966_/B _7966_/C vssd1 vssd1 vccd1 vccd1 _7968_/C sky130_fd_sc_hd__a21o_1
XFILLER_14_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8741__8 vssd1 vssd1 vccd1 vccd1 _8741__8/HI _8836_/A sky130_fd_sc_hd__conb_1
X_6918_ _6918_/A _6918_/B vssd1 vssd1 vccd1 vccd1 _7025_/B sky130_fd_sc_hd__xor2_1
X_7898_ _8206_/A _8335_/A _7897_/C _7897_/D vssd1 vssd1 vccd1 vccd1 _7945_/C sky130_fd_sc_hd__a22o_1
X_6849_ _6857_/A _7432_/A vssd1 vssd1 vccd1 vccd1 _6929_/B sky130_fd_sc_hd__nand2_1
XFILLER_50_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8519_ _7847_/A _8524_/B _7943_/X vssd1 vssd1 vccd1 vccd1 _8520_/B sky130_fd_sc_hd__a21bo_1
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8749__16 vssd1 vssd1 vccd1 vccd1 _8749__16/HI _8844_/A sky130_fd_sc_hd__conb_1
XFILLER_85_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5180_ _5237_/A _5186_/A _5202_/C _5180_/D vssd1 vssd1 vccd1 vccd1 _5180_/X sky130_fd_sc_hd__or4_1
XFILLER_68_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8870_ _8870_/A _4380_/Y vssd1 vssd1 vccd1 vccd1 io_out[7] sky130_fd_sc_hd__ebufn_8
XFILLER_64_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7821_ _7822_/A _7822_/B vssd1 vssd1 vccd1 vccd1 _7934_/A sky130_fd_sc_hd__or2_1
X_8763__30 vssd1 vssd1 vccd1 vccd1 _8763__30/HI _8858_/A sky130_fd_sc_hd__conb_1
XFILLER_91_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4964_ _5107_/A _4964_/B vssd1 vssd1 vccd1 vccd1 _5131_/A sky130_fd_sc_hd__or2_2
X_7752_ _8203_/A _7886_/A vssd1 vssd1 vccd1 vccd1 _7781_/A sky130_fd_sc_hd__nand2_1
X_6703_ _6703_/A _6703_/B vssd1 vssd1 vccd1 vccd1 _6704_/C sky130_fd_sc_hd__xnor2_2
XFILLER_51_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4895_ _4904_/B vssd1 vssd1 vccd1 vccd1 _5047_/B sky130_fd_sc_hd__clkbuf_2
X_7683_ _7683_/A vssd1 vssd1 vccd1 vccd1 _7711_/A sky130_fd_sc_hd__buf_2
X_6634_ _8619_/Q _8702_/Q vssd1 vssd1 vccd1 vccd1 _6635_/B sky130_fd_sc_hd__or2b_1
X_6565_ _6565_/A _7630_/B vssd1 vssd1 vccd1 vccd1 _6588_/B sky130_fd_sc_hd__nand2_1
X_6496_ _6515_/B vssd1 vssd1 vccd1 vccd1 _6526_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_8304_ _8304_/A _8474_/A vssd1 vssd1 vccd1 vccd1 _8304_/Y sky130_fd_sc_hd__nor2_1
X_5516_ _5874_/A _5792_/B _5483_/B _5515_/Y vssd1 vssd1 vccd1 vccd1 _5523_/A sky130_fd_sc_hd__a31o_1
X_8235_ _8235_/A _8235_/B vssd1 vssd1 vccd1 vccd1 _8236_/B sky130_fd_sc_hd__nand2_1
X_5447_ _5447_/A _5447_/B vssd1 vssd1 vccd1 vccd1 _5475_/A sky130_fd_sc_hd__nor2_2
X_8166_ _8365_/B vssd1 vssd1 vccd1 vccd1 _8166_/X sky130_fd_sc_hd__clkbuf_2
X_5378_ _8656_/Q vssd1 vssd1 vccd1 vccd1 _5426_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_101_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7117_ _7116_/B _7117_/B vssd1 vssd1 vccd1 vccd1 _7117_/X sky130_fd_sc_hd__and2b_1
X_8097_ _8106_/B _8097_/B vssd1 vssd1 vccd1 vccd1 _8098_/B sky130_fd_sc_hd__xnor2_1
XFILLER_101_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7048_ _7299_/A _7045_/Y _7046_/X _7047_/X vssd1 vssd1 vccd1 vccd1 _7048_/X sky130_fd_sc_hd__o211a_1
XFILLER_59_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4680_ _8602_/Q vssd1 vssd1 vccd1 vccd1 _5185_/A sky130_fd_sc_hd__inv_2
X_6350_ _6350_/A _6350_/B vssd1 vssd1 vccd1 vccd1 _6350_/Y sky130_fd_sc_hd__nand2_1
X_5301_ _5301_/A _5359_/A _5301_/C vssd1 vssd1 vccd1 vccd1 _5302_/A sky130_fd_sc_hd__and3_1
X_6281_ _6281_/A _6281_/B vssd1 vssd1 vccd1 vccd1 _6282_/B sky130_fd_sc_hd__xnor2_2
XFILLER_5_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5232_ _5227_/C _5230_/X _5231_/X _5214_/A vssd1 vssd1 vccd1 vccd1 _5232_/X sky130_fd_sc_hd__o22a_1
X_8020_ _8020_/A _8020_/B vssd1 vssd1 vccd1 vccd1 _8098_/A sky130_fd_sc_hd__and2_1
X_5163_ _4702_/A _4928_/A _5159_/X _5162_/X vssd1 vssd1 vccd1 vccd1 _5163_/X sky130_fd_sc_hd__o31a_1
XFILLER_68_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5094_ _5220_/A _5245_/B _5092_/X _5093_/X vssd1 vssd1 vccd1 vccd1 _5094_/X sky130_fd_sc_hd__o31a_1
XFILLER_83_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8922_ _8922_/A _4441_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[21] sky130_fd_sc_hd__ebufn_8
X_8853_ _8853_/A _4360_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[22] sky130_fd_sc_hd__ebufn_8
XFILLER_71_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7804_ _7804_/A _7804_/B vssd1 vssd1 vccd1 vccd1 _7805_/A sky130_fd_sc_hd__xor2_1
XFILLER_24_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5996_ _6001_/A vssd1 vssd1 vccd1 vccd1 _6219_/S sky130_fd_sc_hd__dlymetal6s2s_1
X_4947_ _5073_/A _5044_/C vssd1 vssd1 vccd1 vccd1 _4970_/B sky130_fd_sc_hd__or2_1
XFILLER_52_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7735_ _7831_/B _7735_/B vssd1 vssd1 vccd1 vccd1 _7833_/B sky130_fd_sc_hd__nor2_1
XFILLER_20_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7666_ _7722_/A _7666_/B vssd1 vssd1 vccd1 vccd1 _7988_/A sky130_fd_sc_hd__xor2_1
XFILLER_32_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4878_ _4878_/A _4885_/B vssd1 vssd1 vccd1 vccd1 _5126_/A sky130_fd_sc_hd__nor2_1
X_6617_ _6617_/A vssd1 vssd1 vccd1 vccd1 _7443_/A sky130_fd_sc_hd__clkbuf_4
X_7597_ _7597_/A _7597_/B vssd1 vssd1 vccd1 vccd1 _7599_/A sky130_fd_sc_hd__nor2_1
X_6548_ _8709_/Q vssd1 vssd1 vccd1 vccd1 _7516_/A sky130_fd_sc_hd__inv_2
X_6479_ _7520_/A _7514_/A _8709_/Q _7532_/B _7526_/A vssd1 vssd1 vccd1 vccd1 _6479_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_3_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8218_ _8132_/A _8132_/B _8217_/X vssd1 vssd1 vccd1 vccd1 _8223_/A sky130_fd_sc_hd__a21oi_1
XINSDIODE2_0 _5227_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8149_ _8370_/A _8247_/B vssd1 vssd1 vccd1 vccd1 _8152_/A sky130_fd_sc_hd__xnor2_1
XFILLER_87_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5850_ _5850_/A _5850_/B _5690_/C vssd1 vssd1 vccd1 vccd1 _6058_/A sky130_fd_sc_hd__or3b_1
XFILLER_0_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4801_ _6605_/B _4801_/B _4801_/C _4478_/X vssd1 vssd1 vccd1 vccd1 _4802_/A sky130_fd_sc_hd__or4b_1
XFILLER_61_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5781_ _5781_/A _5794_/B vssd1 vssd1 vccd1 vccd1 _5782_/B sky130_fd_sc_hd__xnor2_1
X_7520_ _7520_/A _7526_/B vssd1 vssd1 vccd1 vccd1 _7521_/B sky130_fd_sc_hd__nor2_1
X_4732_ _4478_/X _4733_/S vssd1 vssd1 vccd1 vccd1 _4732_/X sky130_fd_sc_hd__and2b_1
XFILLER_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7451_ _7451_/A _7451_/B vssd1 vssd1 vccd1 vccd1 _7451_/Y sky130_fd_sc_hd__xnor2_1
X_4663_ _5171_/A vssd1 vssd1 vccd1 vccd1 _5226_/B sky130_fd_sc_hd__clkbuf_2
X_6402_ _6402_/A vssd1 vssd1 vccd1 vccd1 _8675_/D sky130_fd_sc_hd__clkbuf_1
X_7382_ _7382_/A _7429_/A _7382_/C vssd1 vssd1 vccd1 vccd1 _7429_/B sky130_fd_sc_hd__nor3_1
X_4594_ _4607_/A vssd1 vssd1 vccd1 vccd1 _4645_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6333_ _6335_/S _6332_/X _6336_/A _6336_/B vssd1 vssd1 vccd1 vccd1 _6333_/X sky130_fd_sc_hd__a211o_1
XFILLER_88_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6264_ _5816_/A _6194_/B _6195_/A vssd1 vssd1 vccd1 vccd1 _6265_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5215_ _5215_/A _5215_/B _5215_/C _5220_/C vssd1 vssd1 vccd1 vccd1 _5215_/X sky130_fd_sc_hd__or4_1
X_8003_ _8022_/A _8003_/B _8003_/C vssd1 vssd1 vccd1 vccd1 _8003_/X sky130_fd_sc_hd__or3_1
XFILLER_69_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6195_ _6195_/A _6195_/B vssd1 vssd1 vccd1 vccd1 _6255_/B sky130_fd_sc_hd__or2_1
X_5146_ _5030_/A _5135_/X _5145_/X vssd1 vssd1 vccd1 vccd1 _5146_/X sky130_fd_sc_hd__o21a_1
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5077_ _5169_/A _5207_/D _5075_/Y _5076_/Y vssd1 vssd1 vccd1 vccd1 _5078_/D sky130_fd_sc_hd__o31a_1
XFILLER_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8905_ _8905_/A _4417_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[4] sky130_fd_sc_hd__ebufn_8
XFILLER_71_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8836_ _8836_/A _4338_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[5] sky130_fd_sc_hd__ebufn_8
XFILLER_25_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5979_ _5979_/A _5979_/B vssd1 vssd1 vccd1 vccd1 _6187_/A sky130_fd_sc_hd__xnor2_1
XFILLER_40_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7718_ _7885_/A _7718_/B vssd1 vssd1 vccd1 vccd1 _7750_/B sky130_fd_sc_hd__xnor2_1
XFILLER_100_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8698_ _8703_/CLK _8698_/D vssd1 vssd1 vccd1 vccd1 _8698_/Q sky130_fd_sc_hd__dfxtp_1
X_7649_ _8515_/A _7649_/B vssd1 vssd1 vccd1 vccd1 _7736_/A sky130_fd_sc_hd__nor2_1
XFILLER_69_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5000_ _5230_/B _5175_/B _5067_/C vssd1 vssd1 vccd1 vccd1 _5227_/D sky130_fd_sc_hd__or3_2
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6951_ _6951_/A _6898_/B vssd1 vssd1 vccd1 vccd1 _6951_/X sky130_fd_sc_hd__or2b_1
XFILLER_93_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6882_ _6882_/A _6882_/B vssd1 vssd1 vccd1 vccd1 _6883_/B sky130_fd_sc_hd__xor2_1
XFILLER_81_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5902_ _5902_/A _5901_/X vssd1 vssd1 vccd1 vccd1 _5903_/B sky130_fd_sc_hd__or2b_1
XFILLER_34_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8621_ _8733_/CLK _8621_/D vssd1 vssd1 vccd1 vccd1 _8621_/Q sky130_fd_sc_hd__dfxtp_2
X_5833_ _5833_/A _6193_/B vssd1 vssd1 vccd1 vccd1 _5833_/Y sky130_fd_sc_hd__nor2_1
XFILLER_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8552_ _7584_/X _8550_/X _8551_/Y vssd1 vssd1 vccd1 vccd1 _8731_/D sky130_fd_sc_hd__o21a_1
X_7503_ _7499_/X _8706_/Q _7497_/X _7502_/X vssd1 vssd1 vccd1 vccd1 _8706_/D sky130_fd_sc_hd__o22a_1
X_5764_ _5763_/A _5841_/A _5763_/C vssd1 vssd1 vccd1 vccd1 _5765_/B sky130_fd_sc_hd__a21oi_1
X_4715_ _4715_/A _4715_/B vssd1 vssd1 vccd1 vccd1 _5149_/S sky130_fd_sc_hd__nand2_2
X_8483_ _8483_/A _8483_/B vssd1 vssd1 vccd1 vccd1 _8484_/B sky130_fd_sc_hd__xnor2_1
X_5695_ _6047_/A _6047_/B _5694_/Y vssd1 vssd1 vccd1 vccd1 _5757_/A sky130_fd_sc_hd__a21boi_2
X_7434_ _7465_/A _7434_/B _7454_/C vssd1 vssd1 vccd1 vccd1 _7434_/X sky130_fd_sc_hd__or3b_1
X_4646_ _4646_/A vssd1 vssd1 vccd1 vccd1 _8600_/D sky130_fd_sc_hd__clkbuf_1
X_7365_ _7454_/B _7364_/C _7364_/B vssd1 vssd1 vccd1 vccd1 _7367_/B sky130_fd_sc_hd__a21o_1
X_4577_ _4577_/A _4577_/B _4577_/C _4577_/D vssd1 vssd1 vccd1 vccd1 _4578_/C sky130_fd_sc_hd__or4_1
X_6316_ _6316_/A _6316_/B vssd1 vssd1 vccd1 vccd1 _6316_/Y sky130_fd_sc_hd__nor2_1
XFILLER_103_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7296_ _7296_/A _7296_/B vssd1 vssd1 vccd1 vccd1 _7484_/B sky130_fd_sc_hd__nor2_1
XFILLER_1_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6247_ _6253_/A _6246_/Y _5981_/B vssd1 vssd1 vccd1 vccd1 _6247_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_97_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6178_ _6178_/A _6178_/B vssd1 vssd1 vccd1 vccd1 _6181_/A sky130_fd_sc_hd__xnor2_1
X_5129_ _5194_/A vssd1 vssd1 vccd1 vccd1 _5237_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_72_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4500_ _5591_/A vssd1 vssd1 vccd1 vccd1 _4808_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5480_ _5480_/A _5480_/B vssd1 vssd1 vccd1 vccd1 _5873_/A sky130_fd_sc_hd__xnor2_4
X_4431_ _4431_/A vssd1 vssd1 vccd1 vccd1 _4431_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4362_ _4363_/A vssd1 vssd1 vccd1 vccd1 _4362_/Y sky130_fd_sc_hd__inv_2
X_7150_ _7141_/A _7141_/C _7141_/B vssd1 vssd1 vccd1 vccd1 _7152_/A sky130_fd_sc_hd__a21boi_1
XFILLER_98_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7081_ _7133_/A _7130_/B vssd1 vssd1 vccd1 vccd1 _7085_/B sky130_fd_sc_hd__xnor2_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6101_ _6101_/A _6101_/B vssd1 vssd1 vccd1 vccd1 _6122_/B sky130_fd_sc_hd__nor2_1
XFILLER_86_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6032_ _5941_/A _5739_/B _5673_/Y vssd1 vssd1 vccd1 vccd1 _6033_/B sky130_fd_sc_hd__a21o_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7983_ _8023_/B _7982_/C _7982_/A vssd1 vssd1 vccd1 vccd1 _8003_/B sky130_fd_sc_hd__a21oi_1
X_6934_ _6934_/A _6934_/B vssd1 vssd1 vccd1 vccd1 _6935_/B sky130_fd_sc_hd__xnor2_1
XFILLER_54_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8604_ _8677_/CLK _8604_/D vssd1 vssd1 vccd1 vccd1 _8604_/Q sky130_fd_sc_hd__dfxtp_1
X_6865_ _6820_/B _6865_/B vssd1 vssd1 vccd1 vccd1 _6865_/X sky130_fd_sc_hd__and2b_1
X_6796_ _7324_/A vssd1 vssd1 vccd1 vccd1 _7102_/B sky130_fd_sc_hd__buf_2
X_5816_ _5816_/A _5816_/B vssd1 vssd1 vccd1 vccd1 _5819_/A sky130_fd_sc_hd__xnor2_2
X_5747_ _5945_/A _5747_/B _5747_/C _5747_/D vssd1 vssd1 vccd1 vccd1 _5838_/A sky130_fd_sc_hd__and4_1
XFILLER_10_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8535_ _8544_/A _8728_/Q vssd1 vssd1 vccd1 vccd1 _8535_/Y sky130_fd_sc_hd__nor2_1
XFILLER_41_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8466_ _8466_/A _8466_/B vssd1 vssd1 vccd1 vccd1 _8467_/B sky130_fd_sc_hd__xnor2_1
X_7417_ _7417_/A _7417_/B vssd1 vssd1 vccd1 vccd1 _7418_/B sky130_fd_sc_hd__xnor2_1
X_5678_ _5678_/A _5678_/B vssd1 vssd1 vccd1 vccd1 _5680_/B sky130_fd_sc_hd__xnor2_1
X_4629_ _8594_/Q _8593_/Q _4623_/B _8595_/Q vssd1 vssd1 vccd1 vccd1 _4630_/C sky130_fd_sc_hd__a31o_1
X_8397_ _8337_/B _8397_/B vssd1 vssd1 vccd1 vccd1 _8404_/B sky130_fd_sc_hd__and2b_1
X_7348_ _7349_/A _7348_/B _7348_/C vssd1 vssd1 vccd1 vccd1 _7355_/B sky130_fd_sc_hd__and3_1
X_7279_ _7279_/A _7279_/B vssd1 vssd1 vccd1 vccd1 _7493_/A sky130_fd_sc_hd__xnor2_1
XFILLER_77_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4980_ _4999_/A vssd1 vssd1 vccd1 vccd1 _5238_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_63_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6650_ _6768_/A _6650_/B vssd1 vssd1 vccd1 vccd1 _6651_/B sky130_fd_sc_hd__nor2_1
X_6581_ _6734_/A _7075_/A vssd1 vssd1 vccd1 vccd1 _6893_/B sky130_fd_sc_hd__nand2_1
X_5601_ _7652_/B _8661_/Q vssd1 vssd1 vccd1 vccd1 _5619_/A sky130_fd_sc_hd__or2b_1
X_5532_ _5532_/A _5532_/B vssd1 vssd1 vccd1 vccd1 _5532_/X sky130_fd_sc_hd__xor2_1
X_8320_ _8223_/A _8223_/B _8319_/Y vssd1 vssd1 vccd1 vccd1 _8326_/A sky130_fd_sc_hd__o21ai_2
X_8251_ _8087_/B _8174_/B _8172_/Y vssd1 vssd1 vccd1 vccd1 _8253_/B sky130_fd_sc_hd__a21o_1
X_5463_ _5480_/A _5480_/B _5450_/A vssd1 vssd1 vccd1 vccd1 _5477_/A sky130_fd_sc_hd__a21o_1
XFILLER_99_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7202_ _7202_/A _7202_/B vssd1 vssd1 vccd1 vccd1 _7475_/A sky130_fd_sc_hd__nor2_1
X_4414_ _4432_/A vssd1 vssd1 vccd1 vccd1 _4419_/A sky130_fd_sc_hd__buf_2
X_8182_ _8187_/A _8187_/B vssd1 vssd1 vccd1 vccd1 _8183_/B sky130_fd_sc_hd__xor2_1
X_5394_ _8657_/Q vssd1 vssd1 vccd1 vccd1 _5615_/A sky130_fd_sc_hd__inv_2
X_4345_ input1/X vssd1 vssd1 vccd1 vccd1 _4370_/A sky130_fd_sc_hd__clkbuf_2
X_7133_ _7133_/A _7254_/C _7133_/C vssd1 vssd1 vccd1 vccd1 _7133_/X sky130_fd_sc_hd__and3_1
XFILLER_98_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7064_ _7432_/B _7261_/B vssd1 vssd1 vccd1 vccd1 _7069_/A sky130_fd_sc_hd__nand2_1
XFILLER_67_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6015_ _6061_/A _6016_/B vssd1 vssd1 vccd1 vccd1 _6312_/A sky130_fd_sc_hd__or2_1
XFILLER_94_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7966_ _8025_/A _7966_/B _7966_/C vssd1 vssd1 vccd1 vccd1 _8025_/B sky130_fd_sc_hd__nand3_1
X_6917_ _6917_/A _6917_/B vssd1 vssd1 vccd1 vccd1 _6918_/B sky130_fd_sc_hd__xnor2_1
X_7897_ _8206_/A _8335_/A _7897_/C _7897_/D vssd1 vssd1 vccd1 vccd1 _7945_/B sky130_fd_sc_hd__nand4_1
X_6848_ _6848_/A _6848_/B vssd1 vssd1 vccd1 vccd1 _7432_/A sky130_fd_sc_hd__nand2_2
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6779_ _6868_/A _6779_/B vssd1 vssd1 vccd1 vccd1 _6869_/A sky130_fd_sc_hd__xnor2_1
X_8518_ _8518_/A _8518_/B vssd1 vssd1 vccd1 vccd1 _8524_/B sky130_fd_sc_hd__xnor2_1
X_8449_ _8321_/A _7878_/A _7761_/Y vssd1 vssd1 vccd1 vccd1 _8450_/C sky130_fd_sc_hd__o21ai_1
XFILLER_2_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7820_ _7661_/X _7748_/Y _7923_/B vssd1 vssd1 vccd1 vccd1 _7822_/B sky130_fd_sc_hd__a21bo_1
X_4963_ _5200_/B _4963_/B vssd1 vssd1 vccd1 vccd1 _5180_/D sky130_fd_sc_hd__or2_1
XFILLER_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7751_ _8118_/A vssd1 vssd1 vccd1 vccd1 _8203_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_24_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6702_ _6682_/X _6702_/B vssd1 vssd1 vccd1 vccd1 _6703_/B sky130_fd_sc_hd__and2b_1
X_7682_ _8605_/Q _8729_/Q vssd1 vssd1 vccd1 vccd1 _7683_/A sky130_fd_sc_hd__or2b_1
X_4894_ _5233_/B _5200_/A vssd1 vssd1 vccd1 vccd1 _4993_/A sky130_fd_sc_hd__or2_1
X_6633_ _8702_/Q _8619_/Q vssd1 vssd1 vccd1 vccd1 _6637_/A sky130_fd_sc_hd__or2b_1
XFILLER_32_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6564_ _6564_/A vssd1 vssd1 vccd1 vccd1 _6588_/A sky130_fd_sc_hd__clkbuf_2
X_6495_ _8697_/Q vssd1 vssd1 vccd1 vccd1 _6515_/B sky130_fd_sc_hd__inv_2
X_8303_ _8460_/A _8303_/B vssd1 vssd1 vccd1 vccd1 _8317_/A sky130_fd_sc_hd__nor2_1
X_5515_ _5566_/A _5784_/A vssd1 vssd1 vccd1 vccd1 _5515_/Y sky130_fd_sc_hd__nor2_1
X_5446_ _8672_/Q _7677_/B vssd1 vssd1 vccd1 vccd1 _5447_/B sky130_fd_sc_hd__and2_1
X_8234_ _8235_/A _8235_/B vssd1 vssd1 vccd1 vccd1 _8345_/B sky130_fd_sc_hd__or2_2
XFILLER_87_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5377_ _6368_/B _5367_/Y _5376_/Y _8558_/A vssd1 vssd1 vccd1 vccd1 _8655_/D sky130_fd_sc_hd__a211o_1
X_8165_ _8080_/A _8080_/B _8081_/A vssd1 vssd1 vccd1 vccd1 _8178_/A sky130_fd_sc_hd__a21oi_1
XFILLER_99_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7116_ _7117_/B _7116_/B vssd1 vssd1 vccd1 vccd1 _7162_/B sky130_fd_sc_hd__xnor2_1
XFILLER_59_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8096_ _8096_/A _8096_/B vssd1 vssd1 vccd1 vccd1 _8097_/B sky130_fd_sc_hd__xnor2_1
X_7047_ _7047_/A _6941_/A vssd1 vssd1 vccd1 vccd1 _7047_/X sky130_fd_sc_hd__or2b_1
XFILLER_86_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7949_ _7881_/B _7881_/C _7881_/A vssd1 vssd1 vccd1 vccd1 _7968_/A sky130_fd_sc_hd__a21bo_1
XFILLER_42_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8809__76 vssd1 vssd1 vccd1 vccd1 _8809__76/HI _8918_/A sky130_fd_sc_hd__conb_1
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5300_ _8635_/Q _8634_/Q vssd1 vssd1 vccd1 vccd1 _5301_/C sky130_fd_sc_hd__nand2_1
X_6280_ _6280_/A _6280_/B vssd1 vssd1 vccd1 vccd1 _6281_/B sky130_fd_sc_hd__xnor2_1
XFILLER_102_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5231_ _5231_/A _5231_/B _5244_/C _5231_/D vssd1 vssd1 vccd1 vccd1 _5231_/X sky130_fd_sc_hd__or4_1
XFILLER_69_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5162_ _5220_/A _5162_/B _5162_/C vssd1 vssd1 vccd1 vccd1 _5162_/X sky130_fd_sc_hd__or3_1
X_5093_ _4942_/A _5208_/A _5084_/X _4958_/B _4665_/A vssd1 vssd1 vccd1 vccd1 _5093_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_96_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8921_ _8921_/A _4440_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[20] sky130_fd_sc_hd__ebufn_8
X_8823__90 vssd1 vssd1 vccd1 vccd1 _8823__90/HI _8932_/A sky130_fd_sc_hd__conb_1
XFILLER_37_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8852_ _8852_/A _4359_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[21] sky130_fd_sc_hd__ebufn_8
XFILLER_37_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7803_ _7741_/A _7738_/X _7741_/B _7739_/A vssd1 vssd1 vccd1 vccd1 _7804_/B sky130_fd_sc_hd__a31o_2
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5995_ _6202_/A _6202_/B vssd1 vssd1 vccd1 vccd1 _6000_/A sky130_fd_sc_hd__xor2_2
X_7734_ _7734_/A _7734_/B vssd1 vssd1 vccd1 vccd1 _7735_/B sky130_fd_sc_hd__and2_1
X_4946_ _5171_/C _5218_/B _5044_/C vssd1 vssd1 vccd1 vccd1 _4946_/X sky130_fd_sc_hd__or3_1
XFILLER_33_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4877_ _5171_/B _4877_/B _5207_/A vssd1 vssd1 vccd1 vccd1 _4996_/A sky130_fd_sc_hd__or3_1
X_7665_ _7835_/A vssd1 vssd1 vccd1 vccd1 _8281_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6616_ _7028_/A _6617_/A vssd1 vssd1 vccd1 vccd1 _6800_/A sky130_fd_sc_hd__nand2_1
XFILLER_20_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7596_ _8717_/Q _7596_/B vssd1 vssd1 vccd1 vccd1 _7597_/B sky130_fd_sc_hd__and2b_1
X_6547_ _8605_/Q _8709_/Q vssd1 vssd1 vccd1 vccd1 _6593_/A sky130_fd_sc_hd__nand2b_2
X_6478_ _8712_/Q vssd1 vssd1 vccd1 vccd1 _7526_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5429_ _5429_/A _5429_/B vssd1 vssd1 vccd1 vccd1 _5429_/X sky130_fd_sc_hd__or2_1
X_8217_ _8217_/A _8331_/A _8410_/B vssd1 vssd1 vccd1 vccd1 _8217_/X sky130_fd_sc_hd__and3_1
X_8148_ _8196_/A _8283_/A _8147_/X vssd1 vssd1 vccd1 vccd1 _8247_/B sky130_fd_sc_hd__o21ba_1
XINSDIODE2_1 _5227_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8079_ _8079_/A _8079_/B vssd1 vssd1 vccd1 vccd1 _8080_/B sky130_fd_sc_hd__or2_1
XFILLER_74_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_0_0_wb_clk_i clkbuf_4_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _8672_/CLK
+ sky130_fd_sc_hd__clkbuf_2
X_4800_ _4692_/A _4687_/B _4718_/A _4697_/X vssd1 vssd1 vccd1 vccd1 _4801_/C sky130_fd_sc_hd__o211a_1
XFILLER_61_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5780_ _5780_/A _5780_/B _5780_/C vssd1 vssd1 vccd1 vccd1 _5794_/B sky130_fd_sc_hd__and3_2
X_4731_ _4729_/X _4730_/Y _4672_/X vssd1 vssd1 vccd1 vccd1 _8610_/D sky130_fd_sc_hd__o21a_1
X_7450_ _7450_/A _7450_/B vssd1 vssd1 vccd1 vccd1 _7451_/B sky130_fd_sc_hd__xnor2_1
X_4662_ _4662_/A _8609_/Q _4480_/C vssd1 vssd1 vccd1 vccd1 _4668_/B sky130_fd_sc_hd__or3b_1
X_6401_ _8675_/Q _6401_/B vssd1 vssd1 vccd1 vccd1 _6402_/A sky130_fd_sc_hd__and2b_1
X_7381_ _7378_/Y _7379_/X _7346_/Y _7347_/X vssd1 vssd1 vccd1 vccd1 _7382_/C sky130_fd_sc_hd__o211a_1
X_4593_ _8584_/Q _4598_/C vssd1 vssd1 vccd1 vccd1 _4597_/A sky130_fd_sc_hd__and2_1
X_6332_ _6332_/A _6332_/B _6332_/C vssd1 vssd1 vccd1 vccd1 _6332_/X sky130_fd_sc_hd__or3_1
X_6263_ _6197_/A _6262_/Y _6198_/B _6198_/A vssd1 vssd1 vccd1 vccd1 _6266_/A sky130_fd_sc_hd__a22oi_1
X_5214_ _5214_/A _5229_/C vssd1 vssd1 vccd1 vccd1 _5220_/C sky130_fd_sc_hd__or2_1
X_8002_ _8084_/A _8002_/B vssd1 vssd1 vccd1 vccd1 _8003_/C sky130_fd_sc_hd__xor2_1
X_6194_ _6194_/A _6194_/B vssd1 vssd1 vccd1 vccd1 _6195_/B sky130_fd_sc_hd__and2_1
X_5145_ _5205_/A _5141_/X _5143_/X _5144_/X _4710_/A vssd1 vssd1 vccd1 vccd1 _5145_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_84_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5076_ _5047_/A _5047_/B _5068_/Y _5175_/A _5226_/B vssd1 vssd1 vccd1 vccd1 _5076_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_56_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8904_ _8904_/A _4419_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[3] sky130_fd_sc_hd__ebufn_8
X_8835_ _8835_/A _4337_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[4] sky130_fd_sc_hd__ebufn_8
XFILLER_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5978_ _5978_/A _5978_/B vssd1 vssd1 vccd1 vccd1 _5979_/B sky130_fd_sc_hd__xor2_1
XFILLER_40_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8697_ _8703_/CLK _8697_/D vssd1 vssd1 vccd1 vccd1 _8697_/Q sky130_fd_sc_hd__dfxtp_1
X_4929_ _4844_/A _4896_/A _5047_/B vssd1 vssd1 vccd1 vccd1 _5073_/A sky130_fd_sc_hd__a21oi_2
X_7717_ _8515_/D _7796_/C _7716_/X vssd1 vssd1 vccd1 vccd1 _7718_/B sky130_fd_sc_hd__o21a_1
XFILLER_100_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7648_ _8066_/A _8063_/A vssd1 vssd1 vccd1 vccd1 _7649_/B sky130_fd_sc_hd__nand2_1
XFILLER_20_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7579_ _7596_/B _7590_/A _8721_/Q vssd1 vssd1 vccd1 vccd1 _7579_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_102_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6950_ _6950_/A _6921_/B vssd1 vssd1 vccd1 vccd1 _6950_/X sky130_fd_sc_hd__or2b_1
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5901_ _5901_/A _5901_/B _5901_/C vssd1 vssd1 vccd1 vccd1 _5901_/X sky130_fd_sc_hd__or3_1
X_6881_ _7349_/A _7083_/B _6879_/Y _6880_/X vssd1 vssd1 vccd1 vccd1 _6882_/B sky130_fd_sc_hd__o211a_1
X_8620_ _8733_/CLK _8620_/D vssd1 vssd1 vccd1 vccd1 _8620_/Q sky130_fd_sc_hd__dfxtp_2
X_5832_ _5944_/B vssd1 vssd1 vccd1 vccd1 _5953_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_61_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5763_ _5763_/A _5841_/A _5763_/C vssd1 vssd1 vccd1 vccd1 _5924_/A sky130_fd_sc_hd__and3_1
X_8551_ _8547_/A _8574_/A _4785_/A vssd1 vssd1 vccd1 vccd1 _8551_/Y sky130_fd_sc_hd__a21oi_1
X_4714_ _4714_/A _5029_/A vssd1 vssd1 vccd1 vccd1 _4715_/B sky130_fd_sc_hd__or2_1
X_7502_ _7510_/A _7505_/B _7502_/C vssd1 vssd1 vccd1 vccd1 _7502_/X sky130_fd_sc_hd__and3_1
X_8482_ _8421_/A _8480_/X _8481_/X vssd1 vssd1 vccd1 vccd1 _8483_/B sky130_fd_sc_hd__o21a_1
X_5694_ _5694_/A _5694_/B vssd1 vssd1 vccd1 vccd1 _5694_/Y sky130_fd_sc_hd__nand2_1
X_7433_ _7431_/Y _7432_/X _7010_/A vssd1 vssd1 vccd1 vccd1 _7460_/A sky130_fd_sc_hd__a21o_1
X_4645_ _4648_/B _4645_/B _4645_/C vssd1 vssd1 vccd1 vccd1 _4646_/A sky130_fd_sc_hd__and3b_1
X_7364_ _7454_/B _7364_/B _7364_/C vssd1 vssd1 vccd1 vccd1 _7447_/C sky130_fd_sc_hd__nand3_1
X_4576_ _8597_/Q _8600_/Q _8599_/Q vssd1 vssd1 vccd1 vccd1 _4577_/D sky130_fd_sc_hd__or3_1
X_6315_ _6315_/A _6320_/A _6320_/B _6320_/C vssd1 vssd1 vccd1 vccd1 _6336_/B sky130_fd_sc_hd__or4_2
X_7295_ _7295_/A _7295_/B _7295_/C vssd1 vssd1 vccd1 vccd1 _7296_/B sky130_fd_sc_hd__and3_1
XFILLER_39_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6246_ _5981_/A _5531_/A _5479_/Y vssd1 vssd1 vccd1 vccd1 _6246_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_69_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6177_ _6177_/A _6268_/B vssd1 vssd1 vccd1 vccd1 _6178_/B sky130_fd_sc_hd__xnor2_1
X_5128_ _5218_/B _5128_/B _5118_/B vssd1 vssd1 vccd1 vccd1 _5128_/X sky130_fd_sc_hd__or3b_1
XFILLER_57_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5059_ _5106_/B _5143_/B vssd1 vssd1 vccd1 vccd1 _5059_/X sky130_fd_sc_hd__or2_1
XFILLER_37_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4430_ _4431_/A vssd1 vssd1 vccd1 vccd1 _4430_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4361_ _4363_/A vssd1 vssd1 vccd1 vccd1 _4361_/Y sky130_fd_sc_hd__inv_2
X_6100_ _6119_/A _6119_/B _6099_/C vssd1 vssd1 vccd1 vccd1 _6101_/B sky130_fd_sc_hd__a21oi_1
X_7080_ _7080_/A vssd1 vssd1 vccd1 vccd1 _7172_/C sky130_fd_sc_hd__clkbuf_2
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6031_ _6097_/B _6096_/B vssd1 vssd1 vccd1 vccd1 _6034_/B sky130_fd_sc_hd__nor2_1
XFILLER_39_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7982_ _7982_/A _8023_/B _7982_/C vssd1 vssd1 vccd1 vccd1 _8022_/A sky130_fd_sc_hd__and3_1
X_6933_ _7027_/A _7027_/B vssd1 vssd1 vccd1 vccd1 _6934_/B sky130_fd_sc_hd__xor2_1
XFILLER_81_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6864_ _7096_/A _6945_/B vssd1 vssd1 vccd1 vccd1 _7115_/B sky130_fd_sc_hd__xor2_1
X_8603_ _8703_/CLK _8603_/D vssd1 vssd1 vccd1 vccd1 _8603_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5815_ _5970_/B _5863_/B vssd1 vssd1 vccd1 vccd1 _5816_/B sky130_fd_sc_hd__xnor2_2
XFILLER_34_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6795_ _6795_/A _6727_/A vssd1 vssd1 vccd1 vccd1 _6924_/A sky130_fd_sc_hd__or2b_1
X_5746_ _5746_/A _5746_/B vssd1 vssd1 vccd1 vccd1 _5747_/D sky130_fd_sc_hd__or2_1
XFILLER_22_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8534_ _7846_/Y _8533_/B _8533_/Y _8525_/A _8525_/B vssd1 vssd1 vccd1 vccd1 _8534_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_41_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8465_ _8465_/A _8465_/B vssd1 vssd1 vccd1 vccd1 _8466_/B sky130_fd_sc_hd__xnor2_1
X_5677_ _6038_/A _6035_/B vssd1 vssd1 vccd1 vccd1 _5680_/A sky130_fd_sc_hd__nor2_1
X_7416_ _7416_/A _7416_/B vssd1 vssd1 vccd1 vccd1 _7417_/B sky130_fd_sc_hd__xor2_1
X_4628_ _8594_/Q _8595_/Q _4628_/C vssd1 vssd1 vccd1 vccd1 _4632_/B sky130_fd_sc_hd__and3_1
X_8396_ _8396_/A _8396_/B vssd1 vssd1 vccd1 vccd1 _8404_/A sky130_fd_sc_hd__and2_1
XFILLER_104_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7347_ _7347_/A _7347_/B _7347_/C _7347_/D vssd1 vssd1 vccd1 vccd1 _7347_/X sky130_fd_sc_hd__or4_1
X_4559_ _8633_/Q _4563_/B vssd1 vssd1 vccd1 vccd1 _4560_/A sky130_fd_sc_hd__and2_1
XFILLER_103_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7278_ _7278_/A _7278_/B vssd1 vssd1 vccd1 vccd1 _7495_/A sky130_fd_sc_hd__xnor2_2
XFILLER_103_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6229_ _6229_/A _6229_/B vssd1 vssd1 vccd1 vccd1 _6230_/B sky130_fd_sc_hd__xnor2_4
XFILLER_85_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8784__51 vssd1 vssd1 vccd1 vccd1 _8784__51/HI _8893_/A sky130_fd_sc_hd__conb_1
XFILLER_82_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6580_ _6670_/A vssd1 vssd1 vccd1 vccd1 _7075_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_31_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5600_ _5660_/A _5661_/A _5661_/B _5599_/X vssd1 vssd1 vccd1 vccd1 _5605_/A sky130_fd_sc_hd__a31o_1
X_5531_ _5531_/A _5781_/A vssd1 vssd1 vccd1 vccd1 _5532_/B sky130_fd_sc_hd__xnor2_1
X_8250_ _8278_/A _8250_/B vssd1 vssd1 vccd1 vccd1 _8253_/A sky130_fd_sc_hd__xor2_1
X_7201_ _7201_/A _7201_/B vssd1 vssd1 vccd1 vccd1 _7202_/B sky130_fd_sc_hd__and2_1
XFILLER_8_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5462_ _5480_/A _5480_/B vssd1 vssd1 vccd1 vccd1 _5874_/B sky130_fd_sc_hd__xor2_4
X_5393_ _6503_/A _5434_/B vssd1 vssd1 vccd1 vccd1 _5398_/A sky130_fd_sc_hd__nor2_2
X_4413_ _4413_/A vssd1 vssd1 vccd1 vccd1 _4413_/Y sky130_fd_sc_hd__inv_2
X_8181_ _8181_/A _8181_/B vssd1 vssd1 vccd1 vccd1 _8187_/B sky130_fd_sc_hd__xnor2_2
X_7132_ _7132_/A vssd1 vssd1 vccd1 vccd1 _7254_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_4344_ _4344_/A vssd1 vssd1 vccd1 vccd1 _4344_/Y sky130_fd_sc_hd__inv_2
X_7063_ _7065_/A _7063_/B vssd1 vssd1 vccd1 vccd1 _7261_/B sky130_fd_sc_hd__nor2_2
XFILLER_100_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6014_ _6160_/A _6014_/B vssd1 vssd1 vccd1 vccd1 _6016_/B sky130_fd_sc_hd__xnor2_1
XFILLER_67_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7965_ _7965_/A _7965_/B vssd1 vssd1 vccd1 vccd1 _7966_/C sky130_fd_sc_hd__xnor2_1
XFILLER_42_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6916_ _6916_/A _6916_/B vssd1 vssd1 vccd1 vccd1 _6917_/B sky130_fd_sc_hd__xor2_1
X_7896_ _7946_/B _7946_/C _7946_/A vssd1 vssd1 vccd1 vccd1 _7897_/D sky130_fd_sc_hd__a21o_1
X_6847_ _7095_/A vssd1 vssd1 vccd1 vccd1 _7039_/A sky130_fd_sc_hd__clkbuf_2
X_6778_ _7004_/A _6884_/A vssd1 vssd1 vccd1 vccd1 _6779_/B sky130_fd_sc_hd__xnor2_2
Xclkbuf_4_13_0_wb_clk_i clkbuf_3_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8703_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_52_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5729_ _5729_/A _5729_/B vssd1 vssd1 vccd1 vccd1 _5751_/A sky130_fd_sc_hd__nand2_1
X_8517_ _8525_/A _8525_/B _8523_/B vssd1 vssd1 vccd1 vccd1 _8517_/X sky130_fd_sc_hd__or3_1
X_8448_ _8448_/A _8448_/B vssd1 vssd1 vccd1 vccd1 _8452_/A sky130_fd_sc_hd__xnor2_1
X_8379_ _8439_/B _8379_/B vssd1 vssd1 vccd1 vccd1 _8382_/A sky130_fd_sc_hd__xnor2_1
XFILLER_2_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4962_ _5223_/B vssd1 vssd1 vccd1 vccd1 _5200_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_51_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7750_ _7750_/A _7750_/B vssd1 vssd1 vccd1 vccd1 _7826_/A sky130_fd_sc_hd__or2_1
X_6701_ _7169_/A _7083_/B vssd1 vssd1 vccd1 vccd1 _6703_/A sky130_fd_sc_hd__nand2_1
X_4893_ _4950_/B _4969_/B vssd1 vssd1 vccd1 vccd1 _5200_/A sky130_fd_sc_hd__nand2_2
X_7681_ _7681_/A _7681_/B vssd1 vssd1 vccd1 vccd1 _7712_/A sky130_fd_sc_hd__nor2_2
X_6632_ _6579_/A _6579_/B _6631_/Y vssd1 vssd1 vccd1 vccd1 _6652_/B sky130_fd_sc_hd__a21o_1
XFILLER_20_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6563_ _8615_/Q _8698_/Q vssd1 vssd1 vccd1 vccd1 _6564_/A sky130_fd_sc_hd__or2b_1
X_6494_ _8703_/Q vssd1 vssd1 vccd1 vccd1 _6536_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_8302_ _8390_/A vssd1 vssd1 vccd1 vccd1 _8460_/A sky130_fd_sc_hd__inv_2
X_5514_ _5500_/A _5500_/B _5513_/Y vssd1 vssd1 vccd1 vccd1 _5535_/A sky130_fd_sc_hd__a21bo_1
X_8233_ _8328_/A _8328_/B vssd1 vssd1 vccd1 vccd1 _8235_/B sky130_fd_sc_hd__xnor2_1
X_5445_ _8672_/Q _6603_/B vssd1 vssd1 vccd1 vccd1 _5447_/A sky130_fd_sc_hd__nor2_1
X_8164_ _8190_/A _8164_/B vssd1 vssd1 vccd1 vccd1 _8181_/A sky130_fd_sc_hd__xnor2_2
XFILLER_99_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7115_ _7115_/A _7115_/B vssd1 vssd1 vccd1 vccd1 _7116_/B sky130_fd_sc_hd__xnor2_1
X_5376_ _5372_/X _5374_/X _8673_/Q _6360_/A vssd1 vssd1 vccd1 vccd1 _5376_/Y sky130_fd_sc_hd__a211oi_1
XFILLER_87_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8095_ _8186_/A _8095_/B vssd1 vssd1 vccd1 vccd1 _8096_/B sky130_fd_sc_hd__and2_1
X_7046_ _7046_/A _6940_/A vssd1 vssd1 vccd1 vccd1 _7046_/X sky130_fd_sc_hd__or2b_1
XFILLER_47_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7948_ _7893_/B _7893_/C _7893_/A vssd1 vssd1 vccd1 vccd1 _7978_/A sky130_fd_sc_hd__a21bo_1
XFILLER_27_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8754__21 vssd1 vssd1 vccd1 vccd1 _8754__21/HI _8849_/A sky130_fd_sc_hd__conb_1
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7879_ _8217_/A _7963_/A _7878_/Y vssd1 vssd1 vccd1 vccd1 _7880_/B sky130_fd_sc_hd__a21oi_1
XFILLER_10_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5230_ _5230_/A _5230_/B _5236_/C _5230_/D vssd1 vssd1 vccd1 vccd1 _5230_/X sky130_fd_sc_hd__or4_1
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5161_ _4914_/A _5231_/A _5106_/C _5160_/X _5227_/C vssd1 vssd1 vccd1 vccd1 _5162_/C
+ sky130_fd_sc_hd__o32a_1
XFILLER_69_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5092_ _5173_/A _5106_/B _5238_/B _5106_/C _5200_/C vssd1 vssd1 vccd1 vccd1 _5092_/X
+ sky130_fd_sc_hd__o41a_1
XFILLER_68_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8920_ _8920_/A _4439_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[19] sky130_fd_sc_hd__ebufn_8
X_8851_ _8851_/A _4357_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[20] sky130_fd_sc_hd__ebufn_8
XFILLER_64_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7802_ _8051_/A _7802_/B vssd1 vssd1 vccd1 vccd1 _7804_/A sky130_fd_sc_hd__and2_1
XFILLER_24_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5994_ _6218_/B _5994_/B vssd1 vssd1 vccd1 vccd1 _6202_/B sky130_fd_sc_hd__xor2_1
XFILLER_37_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4945_ _5002_/B vssd1 vssd1 vccd1 vccd1 _5218_/B sky130_fd_sc_hd__buf_2
XFILLER_24_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7733_ _7734_/A _7734_/B vssd1 vssd1 vccd1 vccd1 _7831_/B sky130_fd_sc_hd__nor2_1
XFILLER_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7664_ _7834_/A vssd1 vssd1 vccd1 vccd1 _7835_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4876_ _4876_/A _4904_/A vssd1 vssd1 vccd1 vccd1 _5207_/A sky130_fd_sc_hd__nor2_1
X_6615_ _6835_/A vssd1 vssd1 vccd1 vccd1 _7028_/A sky130_fd_sc_hd__inv_2
X_7595_ _7595_/A vssd1 vssd1 vccd1 vccd1 _8719_/D sky130_fd_sc_hd__clkbuf_1
X_6546_ _6546_/A vssd1 vssd1 vccd1 vccd1 _8704_/D sky130_fd_sc_hd__clkbuf_1
X_6477_ _8710_/Q vssd1 vssd1 vccd1 vccd1 _7514_/A sky130_fd_sc_hd__clkbuf_2
X_5428_ _5427_/A _5433_/S _5427_/C _5432_/B vssd1 vssd1 vccd1 vccd1 _5429_/B sky130_fd_sc_hd__a22oi_1
X_8216_ _8220_/B vssd1 vssd1 vccd1 vccd1 _8410_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_99_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5359_ _5359_/A _5359_/B _5359_/C vssd1 vssd1 vccd1 vccd1 _5360_/A sky130_fd_sc_hd__and3_1
XFILLER_87_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8147_ _8150_/A _7805_/A _8057_/A _7661_/A vssd1 vssd1 vccd1 vccd1 _8147_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_101_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_2 _4464_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8078_ _8078_/A _8078_/B vssd1 vssd1 vccd1 vccd1 _8080_/A sky130_fd_sc_hd__nand2_1
XFILLER_101_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7029_ _7280_/B _6916_/B _6917_/A _6917_/B vssd1 vssd1 vccd1 vccd1 _7317_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_43_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4730_ _4733_/S _4730_/B vssd1 vssd1 vccd1 vccd1 _4730_/Y sky130_fd_sc_hd__nor2_1
XFILLER_14_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4661_ _4661_/A _4763_/A vssd1 vssd1 vccd1 vccd1 _4702_/B sky130_fd_sc_hd__nand2_1
XFILLER_9_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7380_ _7346_/Y _7347_/X _7378_/Y _7379_/X vssd1 vssd1 vccd1 vccd1 _7429_/A sky130_fd_sc_hd__a211oi_2
X_6400_ _6464_/B vssd1 vssd1 vccd1 vccd1 _6401_/B sky130_fd_sc_hd__clkbuf_2
X_6331_ _6331_/A _6332_/A vssd1 vssd1 vccd1 vccd1 _6335_/S sky130_fd_sc_hd__or2b_1
X_4592_ _4592_/A vssd1 vssd1 vccd1 vccd1 _8583_/D sky130_fd_sc_hd__clkbuf_1
X_6262_ _6262_/A vssd1 vssd1 vccd1 vccd1 _6262_/Y sky130_fd_sc_hd__inv_2
X_5213_ _5120_/B _5170_/B _5212_/X _4923_/X vssd1 vssd1 vccd1 vccd1 _5215_/C sky130_fd_sc_hd__o31a_1
X_6193_ _6193_/A _6193_/B vssd1 vssd1 vccd1 vccd1 _6195_/A sky130_fd_sc_hd__nor2_1
X_8001_ _7922_/A _7922_/B _8000_/Y vssd1 vssd1 vccd1 vccd1 _8002_/B sky130_fd_sc_hd__o21ai_1
X_5144_ _5164_/C _5132_/X _5127_/X _4522_/A _5053_/A vssd1 vssd1 vccd1 vccd1 _5144_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_96_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5075_ _5173_/A _4827_/A _4942_/A vssd1 vssd1 vccd1 vccd1 _5075_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_84_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8903_ _8903_/A _4422_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[2] sky130_fd_sc_hd__ebufn_8
X_8834_ _8834_/A _4336_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[3] sky130_fd_sc_hd__ebufn_8
XFILLER_25_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5977_ _6255_/A _6190_/B vssd1 vssd1 vccd1 vccd1 _5978_/B sky130_fd_sc_hd__xnor2_1
X_8696_ _8715_/CLK _8696_/D vssd1 vssd1 vccd1 vccd1 _8696_/Q sky130_fd_sc_hd__dfxtp_1
X_4928_ _4928_/A _5166_/B _4928_/C vssd1 vssd1 vccd1 vccd1 _4928_/X sky130_fd_sc_hd__or3_1
XFILLER_52_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7716_ _8139_/A _8399_/B vssd1 vssd1 vccd1 vccd1 _7716_/X sky130_fd_sc_hd__or2_1
XFILLER_20_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7647_ _8065_/A vssd1 vssd1 vccd1 vccd1 _8063_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_60_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4859_ _4859_/A _4899_/B vssd1 vssd1 vccd1 vccd1 _4864_/B sky130_fd_sc_hd__nor2_1
X_7578_ _7618_/A _7574_/Y _7613_/A _7577_/X vssd1 vssd1 vccd1 vccd1 _7578_/Y sky130_fd_sc_hd__a31oi_1
X_6529_ _6528_/A _6534_/A _6528_/C vssd1 vssd1 vccd1 vccd1 _6529_/X sky130_fd_sc_hd__a21o_1
XFILLER_79_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5900_ _5901_/A _5901_/B _5901_/C vssd1 vssd1 vccd1 vccd1 _5902_/A sky130_fd_sc_hd__o21a_1
X_6880_ _7348_/B vssd1 vssd1 vccd1 vccd1 _6880_/X sky130_fd_sc_hd__clkbuf_2
X_5831_ _6030_/A vssd1 vssd1 vccd1 vccd1 _5831_/X sky130_fd_sc_hd__buf_2
XFILLER_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5762_ _5729_/B _5747_/B _5970_/A vssd1 vssd1 vccd1 vccd1 _5763_/C sky130_fd_sc_hd__o21a_1
XFILLER_22_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8550_ _8550_/A _8550_/B vssd1 vssd1 vccd1 vccd1 _8550_/X sky130_fd_sc_hd__xor2_1
X_4713_ _4714_/A _5029_/A vssd1 vssd1 vccd1 vccd1 _4715_/A sky130_fd_sc_hd__nand2_1
X_7501_ _7501_/A _7501_/B vssd1 vssd1 vccd1 vccd1 _7502_/C sky130_fd_sc_hd__or2_1
X_5693_ _5769_/A _5693_/B vssd1 vssd1 vccd1 vccd1 _6047_/B sky130_fd_sc_hd__nor2_1
X_8481_ _8481_/A _8420_/B vssd1 vssd1 vccd1 vccd1 _8481_/X sky130_fd_sc_hd__or2b_1
X_7432_ _7432_/A _7432_/B _7432_/C vssd1 vssd1 vccd1 vccd1 _7432_/X sky130_fd_sc_hd__or3_1
X_4644_ _8599_/Q _4643_/C _8600_/Q vssd1 vssd1 vccd1 vccd1 _4645_/C sky130_fd_sc_hd__a21o_1
X_7363_ _7362_/A _7362_/B _7362_/C vssd1 vssd1 vccd1 vccd1 _7378_/B sky130_fd_sc_hd__a21oi_1
X_4575_ _8596_/Q _8595_/Q _8598_/Q _8601_/Q vssd1 vssd1 vccd1 vccd1 _4577_/C sky130_fd_sc_hd__or4b_1
X_7294_ _7295_/B _7295_/C _7295_/A vssd1 vssd1 vccd1 vccd1 _7296_/A sky130_fd_sc_hd__a21oi_1
X_6314_ _6305_/A _6305_/B _6306_/X _6309_/Y _6313_/X vssd1 vssd1 vccd1 vccd1 _6320_/C
+ sky130_fd_sc_hd__a2111o_1
XFILLER_89_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6245_ _6245_/A _6245_/B vssd1 vssd1 vccd1 vccd1 _6249_/A sky130_fd_sc_hd__xnor2_1
XFILLER_103_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6176_ _6176_/A _6176_/B vssd1 vssd1 vccd1 vccd1 _6268_/B sky130_fd_sc_hd__xor2_1
XFILLER_84_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5127_ _5127_/A _5220_/B _5212_/B _5127_/D vssd1 vssd1 vccd1 vccd1 _5127_/X sky130_fd_sc_hd__or4_1
XFILLER_69_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5058_ _5086_/B _5078_/C _5155_/A vssd1 vssd1 vccd1 vccd1 _5058_/X sky130_fd_sc_hd__o21a_1
XFILLER_84_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8679_ _8695_/CLK _8679_/D vssd1 vssd1 vccd1 vccd1 _8679_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4360_ _4363_/A vssd1 vssd1 vccd1 vccd1 _4360_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6030_ _6030_/A _6030_/B _6095_/A vssd1 vssd1 vccd1 vccd1 _6096_/B sky130_fd_sc_hd__and3_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7981_ _8023_/A _7980_/C _7980_/A vssd1 vssd1 vccd1 vccd1 _7982_/C sky130_fd_sc_hd__a21o_1
X_6932_ _6932_/A _6932_/B vssd1 vssd1 vccd1 vccd1 _7027_/B sky130_fd_sc_hd__xnor2_1
XFILLER_81_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6863_ _6863_/A _6863_/B vssd1 vssd1 vccd1 vccd1 _6945_/B sky130_fd_sc_hd__xnor2_1
X_8602_ _8703_/CLK _8602_/D vssd1 vssd1 vccd1 vccd1 _8602_/Q sky130_fd_sc_hd__dfxtp_1
X_5814_ _5814_/A vssd1 vssd1 vccd1 vccd1 _5863_/B sky130_fd_sc_hd__clkbuf_2
X_6794_ _6763_/A _6791_/X _6792_/Y _6793_/X vssd1 vssd1 vccd1 vccd1 _6818_/A sky130_fd_sc_hd__a31o_1
XFILLER_22_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5745_ _5820_/A _5745_/B vssd1 vssd1 vccd1 vccd1 _5747_/C sky130_fd_sc_hd__xnor2_1
X_8533_ _8533_/A _8533_/B vssd1 vssd1 vccd1 vccd1 _8533_/Y sky130_fd_sc_hd__nor2_1
X_8464_ _8464_/A _8464_/B vssd1 vssd1 vccd1 vccd1 _8465_/B sky130_fd_sc_hd__xnor2_1
X_5676_ _5682_/A _5676_/B vssd1 vssd1 vccd1 vccd1 _6035_/B sky130_fd_sc_hd__xnor2_1
X_7415_ _7146_/A _7430_/B _7065_/X _7409_/B _7010_/A vssd1 vssd1 vccd1 vccd1 _7416_/B
+ sky130_fd_sc_hd__a221o_1
X_4627_ _8594_/Q _4628_/C _4626_/Y vssd1 vssd1 vccd1 vccd1 _8594_/D sky130_fd_sc_hd__a21oi_1
X_8395_ _8347_/A _8347_/B _8346_/A vssd1 vssd1 vccd1 vccd1 _8481_/A sky130_fd_sc_hd__a21oi_2
X_7346_ _7347_/C vssd1 vssd1 vccd1 vccd1 _7346_/Y sky130_fd_sc_hd__inv_2
XFILLER_89_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4558_ _4558_/A vssd1 vssd1 vccd1 vccd1 _8886_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_104_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7277_ _7279_/A _7279_/B _7276_/X vssd1 vssd1 vccd1 vccd1 _7278_/B sky130_fd_sc_hd__a21oi_2
X_4489_ _4847_/A vssd1 vssd1 vccd1 vccd1 _4749_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6228_ _6278_/A _6278_/B vssd1 vssd1 vccd1 vccd1 _6229_/B sky130_fd_sc_hd__xor2_2
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6159_ _6062_/Y _6306_/A _6306_/B _6158_/X vssd1 vssd1 vccd1 vccd1 _6302_/B sky130_fd_sc_hd__a31o_1
XFILLER_85_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5530_ _5530_/A vssd1 vssd1 vccd1 vccd1 _5781_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_8_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5461_ _6071_/A _5872_/A vssd1 vssd1 vccd1 vccd1 _5501_/A sky130_fd_sc_hd__nand2_1
X_7200_ _7201_/A _7201_/B vssd1 vssd1 vccd1 vccd1 _7202_/A sky130_fd_sc_hd__nor2_1
X_4412_ _4413_/A vssd1 vssd1 vccd1 vccd1 _4412_/Y sky130_fd_sc_hd__inv_2
X_8180_ _8180_/A _8180_/B vssd1 vssd1 vccd1 vccd1 _8181_/B sky130_fd_sc_hd__xor2_2
X_5392_ _7614_/A _5410_/A vssd1 vssd1 vccd1 vccd1 _5397_/A sky130_fd_sc_hd__nor2_1
X_7131_ _7131_/A _7133_/C vssd1 vssd1 vccd1 vccd1 _7173_/B sky130_fd_sc_hd__xnor2_1
X_4343_ _4344_/A vssd1 vssd1 vccd1 vccd1 _4343_/Y sky130_fd_sc_hd__inv_2
X_7062_ _7068_/A _7270_/A vssd1 vssd1 vccd1 vccd1 _7147_/B sky130_fd_sc_hd__nor2_1
XFILLER_59_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6013_ _6013_/A _6013_/B vssd1 vssd1 vccd1 vccd1 _6014_/B sky130_fd_sc_hd__xor2_1
XFILLER_86_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7964_ _8399_/A _8044_/A _7963_/X vssd1 vssd1 vccd1 vccd1 _7965_/B sky130_fd_sc_hd__a21oi_1
XFILLER_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6915_ _7033_/A _6915_/B vssd1 vssd1 vccd1 vccd1 _6917_/A sky130_fd_sc_hd__nor2_1
XFILLER_82_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7895_ _7946_/A _7946_/B _7946_/C vssd1 vssd1 vccd1 vccd1 _7897_/C sky130_fd_sc_hd__nand3_1
X_6846_ _6765_/A _6765_/B _6845_/X vssd1 vssd1 vccd1 vccd1 _6863_/A sky130_fd_sc_hd__a21o_1
XFILLER_50_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6777_ _7364_/B _7443_/B vssd1 vssd1 vccd1 vccd1 _6884_/A sky130_fd_sc_hd__xnor2_1
X_5728_ _5728_/A _5728_/B vssd1 vssd1 vccd1 vccd1 _5754_/A sky130_fd_sc_hd__nand2_1
X_8516_ _8518_/A _8514_/X _8515_/X vssd1 vssd1 vccd1 vccd1 _8523_/B sky130_fd_sc_hd__a21oi_1
X_5659_ _8660_/Q _4861_/B vssd1 vssd1 vccd1 vccd1 _5660_/B sky130_fd_sc_hd__or2b_1
X_8447_ _8330_/A _8410_/Y _7963_/X vssd1 vssd1 vccd1 vccd1 _8448_/B sky130_fd_sc_hd__o21ba_1
X_8378_ _8378_/A _8378_/B vssd1 vssd1 vccd1 vccd1 _8379_/B sky130_fd_sc_hd__xnor2_1
XFILLER_104_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7329_ _7444_/A _7329_/B vssd1 vssd1 vccd1 vccd1 _7329_/X sky130_fd_sc_hd__and2_1
XFILLER_2_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4961_ _5107_/A _5222_/B vssd1 vssd1 vccd1 vccd1 _5188_/C sky130_fd_sc_hd__or2_1
XFILLER_17_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6700_ _6700_/A vssd1 vssd1 vccd1 vccd1 _7083_/B sky130_fd_sc_hd__buf_2
X_4892_ _4990_/A _4948_/B vssd1 vssd1 vccd1 vccd1 _4969_/B sky130_fd_sc_hd__or2_1
X_7680_ _8607_/Q _8731_/Q vssd1 vssd1 vccd1 vccd1 _7681_/B sky130_fd_sc_hd__and2b_1
X_6631_ _6631_/A _6659_/B vssd1 vssd1 vccd1 vccd1 _6631_/Y sky130_fd_sc_hd__nand2_1
X_6562_ _7065_/A _7335_/A vssd1 vssd1 vccd1 vccd1 _6587_/A sky130_fd_sc_hd__or2_1
X_8301_ _8240_/A _8240_/B _8300_/X vssd1 vssd1 vccd1 vccd1 _8350_/A sky130_fd_sc_hd__a21oi_1
X_6493_ _6498_/A _6500_/A _6491_/Y _6536_/B vssd1 vssd1 vccd1 vccd1 _6493_/X sky130_fd_sc_hd__a31o_1
X_5513_ _5788_/A _5513_/B vssd1 vssd1 vccd1 vccd1 _5513_/Y sky130_fd_sc_hd__nand2_1
X_5444_ _6020_/A vssd1 vssd1 vccd1 vccd1 _6071_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_8232_ _8341_/B _8232_/B vssd1 vssd1 vccd1 vccd1 _8328_/B sky130_fd_sc_hd__nand2_1
X_8163_ _8163_/A _8163_/B vssd1 vssd1 vccd1 vccd1 _8164_/B sky130_fd_sc_hd__xor2_2
X_7114_ _7156_/A _7156_/B _7113_/Y vssd1 vssd1 vccd1 vccd1 _7117_/B sky130_fd_sc_hd__a21o_1
X_5375_ _8672_/Q vssd1 vssd1 vccd1 vccd1 _6360_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_101_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8094_ _8094_/A _8094_/B vssd1 vssd1 vccd1 vccd1 _8095_/B sky130_fd_sc_hd__nand2_1
X_7045_ _7042_/X _7043_/Y _6948_/X _6949_/Y vssd1 vssd1 vccd1 vccd1 _7045_/Y sky130_fd_sc_hd__a211oi_2
XFILLER_86_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7947_ _8206_/A _8335_/A _7897_/D _7946_/X vssd1 vssd1 vccd1 vccd1 _7982_/A sky130_fd_sc_hd__a31o_1
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7878_ _7878_/A _7888_/A vssd1 vssd1 vccd1 vccd1 _7878_/Y sky130_fd_sc_hd__nor2_1
XFILLER_35_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6829_ _6829_/A _6839_/B vssd1 vssd1 vccd1 vccd1 _6931_/B sky130_fd_sc_hd__or2_1
XFILLER_11_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5160_ _5194_/A _5188_/B _5223_/A _5186_/C vssd1 vssd1 vccd1 vccd1 _5160_/X sky130_fd_sc_hd__or4_1
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5091_ _5248_/A _5215_/B _5091_/C vssd1 vssd1 vccd1 vccd1 _5091_/X sky130_fd_sc_hd__or3_1
XFILLER_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8850_ _8850_/A _4356_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[19] sky130_fd_sc_hd__ebufn_8
XFILLER_76_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7801_ _8621_/Q _7577_/X vssd1 vssd1 vccd1 vccd1 _7802_/B sky130_fd_sc_hd__or2b_1
X_5993_ _5993_/A _6001_/A vssd1 vssd1 vccd1 vccd1 _5994_/B sky130_fd_sc_hd__xor2_1
X_4944_ _5222_/A _4979_/A vssd1 vssd1 vccd1 vccd1 _4965_/B sky130_fd_sc_hd__or2_1
XFILLER_52_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7732_ _8139_/A _7796_/C _7841_/A _7841_/B vssd1 vssd1 vccd1 vccd1 _7734_/B sky130_fd_sc_hd__o22a_1
X_7663_ _7725_/A vssd1 vssd1 vccd1 vccd1 _7663_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_32_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4875_ _4919_/A _4937_/B vssd1 vssd1 vccd1 vccd1 _5171_/B sky130_fd_sc_hd__nor2_1
X_6614_ _6614_/A _6744_/A vssd1 vssd1 vccd1 vccd1 _6759_/A sky130_fd_sc_hd__or2_2
X_7594_ _8544_/A _7594_/B vssd1 vssd1 vccd1 vccd1 _7595_/A sky130_fd_sc_hd__and2_1
X_6545_ _7550_/A _6545_/B _6545_/C vssd1 vssd1 vccd1 vccd1 _6546_/A sky130_fd_sc_hd__and3_1
XFILLER_20_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6476_ _8711_/Q vssd1 vssd1 vccd1 vccd1 _7520_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_3_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8215_ _7775_/A _7768_/B _7775_/B _7876_/X _8203_/A vssd1 vssd1 vccd1 vccd1 _8220_/B
+ sky130_fd_sc_hd__o311a_2
X_5427_ _5427_/A _5433_/S _5427_/C _5432_/B vssd1 vssd1 vccd1 vccd1 _5429_/A sky130_fd_sc_hd__and4_1
X_5358_ _8652_/Q _5358_/B vssd1 vssd1 vccd1 vccd1 _5359_/C sky130_fd_sc_hd__nand2_1
XFILLER_87_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8146_ _8150_/A _8146_/B vssd1 vssd1 vccd1 vccd1 _8283_/A sky130_fd_sc_hd__nand2_1
XFILLER_87_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_3 _4464_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8077_ _8161_/A _8077_/B vssd1 vssd1 vccd1 vccd1 _8081_/A sky130_fd_sc_hd__or2_1
X_5289_ _8637_/Q _8636_/Q _5301_/A _6466_/B _8639_/Q vssd1 vssd1 vccd1 vccd1 _5289_/X
+ sky130_fd_sc_hd__a311o_1
X_7028_ _7028_/A vssd1 vssd1 vccd1 vccd1 _7280_/B sky130_fd_sc_hd__buf_2
XFILLER_87_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8814__81 vssd1 vssd1 vccd1 vccd1 _8814__81/HI _8923_/A sky130_fd_sc_hd__conb_1
XFILLER_74_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4660_ _4660_/A _4660_/B _5047_/A _5634_/B vssd1 vssd1 vccd1 vccd1 _4763_/A sky130_fd_sc_hd__or4b_4
XFILLER_80_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6330_ _6324_/X _6329_/X _6325_/X _8665_/Q vssd1 vssd1 vccd1 vccd1 _8665_/D sky130_fd_sc_hd__o2bb2a_1
X_4591_ _4598_/C _4612_/B _4591_/C vssd1 vssd1 vccd1 vccd1 _4592_/A sky130_fd_sc_hd__and3b_1
X_6261_ _6261_/A _6261_/B vssd1 vssd1 vccd1 vccd1 _6267_/A sky130_fd_sc_hd__xnor2_1
X_5212_ _5212_/A _5212_/B vssd1 vssd1 vccd1 vccd1 _5212_/X sky130_fd_sc_hd__or2_1
XFILLER_69_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6192_ _5989_/A _5989_/B _6191_/Y vssd1 vssd1 vccd1 vccd1 _6197_/A sky130_fd_sc_hd__a21bo_1
X_8000_ _8000_/A _8000_/B vssd1 vssd1 vccd1 vccd1 _8000_/Y sky130_fd_sc_hd__nand2_1
X_5143_ _5143_/A _5143_/B _5143_/C vssd1 vssd1 vccd1 vccd1 _5143_/X sky130_fd_sc_hd__or3_1
XFILLER_84_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5074_ _5194_/A vssd1 vssd1 vccd1 vccd1 _5173_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_69_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8902_ _8902_/A _4424_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[1] sky130_fd_sc_hd__ebufn_8
XFILLER_71_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8833_ _8833_/A _4335_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[2] sky130_fd_sc_hd__ebufn_8
XFILLER_52_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5976_ _5976_/A _5976_/B vssd1 vssd1 vccd1 vccd1 _6190_/B sky130_fd_sc_hd__xnor2_2
XFILLER_100_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8695_ _8695_/CLK _8695_/D vssd1 vssd1 vccd1 vccd1 _8695_/Q sky130_fd_sc_hd__dfxtp_1
X_4927_ _5111_/A _5210_/B _4927_/C _4927_/D vssd1 vssd1 vccd1 vccd1 _4928_/C sky130_fd_sc_hd__or4_1
XFILLER_40_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7715_ _8122_/C _8122_/B vssd1 vssd1 vccd1 vccd1 _8399_/B sky130_fd_sc_hd__nand2_1
X_4858_ _5037_/A _5120_/B vssd1 vssd1 vccd1 vccd1 _4991_/B sky130_fd_sc_hd__or2_1
X_7646_ _7656_/A _7656_/B vssd1 vssd1 vccd1 vccd1 _8065_/A sky130_fd_sc_hd__xnor2_2
X_4789_ _8558_/A _4789_/B vssd1 vssd1 vccd1 vccd1 _8621_/D sky130_fd_sc_hd__nor2_1
X_7577_ _8724_/Q vssd1 vssd1 vccd1 vccd1 _7577_/X sky130_fd_sc_hd__clkbuf_2
X_6528_ _6528_/A _6534_/A _6528_/C vssd1 vssd1 vccd1 vccd1 _6541_/A sky130_fd_sc_hd__nand3_1
X_6459_ _8693_/Q _6459_/B vssd1 vssd1 vccd1 vccd1 _6461_/A sky130_fd_sc_hd__and2_1
XFILLER_69_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8129_ _8321_/A _8204_/A vssd1 vssd1 vccd1 vccd1 _8132_/A sky130_fd_sc_hd__nor2_1
XFILLER_87_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5830_ _5830_/A _5854_/B vssd1 vssd1 vccd1 vccd1 _5848_/A sky130_fd_sc_hd__xnor2_1
XFILLER_61_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5761_ _5944_/A vssd1 vssd1 vccd1 vccd1 _5970_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_34_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4712_ _4480_/C _4716_/A _4711_/X _4672_/X vssd1 vssd1 vccd1 vccd1 _8606_/D sky130_fd_sc_hd__o211a_1
X_7500_ _7501_/A _7501_/B vssd1 vssd1 vccd1 vccd1 _7505_/B sky130_fd_sc_hd__nand2_1
X_8480_ _8420_/B _8481_/A vssd1 vssd1 vccd1 vccd1 _8480_/X sky130_fd_sc_hd__and2b_1
X_7431_ _7432_/B _7432_/C _7432_/A vssd1 vssd1 vccd1 vccd1 _7431_/Y sky130_fd_sc_hd__o21ai_1
X_5692_ _5850_/A _5692_/B _5692_/C vssd1 vssd1 vccd1 vccd1 _5693_/B sky130_fd_sc_hd__and3_1
XFILLER_30_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4643_ _8600_/Q _8599_/Q _4643_/C vssd1 vssd1 vccd1 vccd1 _4648_/B sky130_fd_sc_hd__and3_1
X_7362_ _7362_/A _7362_/B _7362_/C vssd1 vssd1 vccd1 vccd1 _7378_/A sky130_fd_sc_hd__and3_1
X_4574_ _8588_/Q _8587_/Q _8590_/Q _8589_/Q vssd1 vssd1 vccd1 vccd1 _4577_/B sky130_fd_sc_hd__or4_1
X_7293_ _7293_/A _7293_/B vssd1 vssd1 vccd1 vccd1 _7295_/A sky130_fd_sc_hd__xnor2_1
X_6313_ _6309_/A _6309_/B _6310_/X _6311_/Y _6312_/X vssd1 vssd1 vccd1 vccd1 _6313_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_89_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6244_ _5992_/A _6218_/Y _5569_/X vssd1 vssd1 vccd1 vccd1 _6245_/B sky130_fd_sc_hd__o21bai_1
XFILLER_69_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6175_ _6175_/A _6270_/B vssd1 vssd1 vccd1 vccd1 _6176_/B sky130_fd_sc_hd__xnor2_1
X_5126_ _5126_/A _5126_/B _5210_/B vssd1 vssd1 vccd1 vccd1 _5127_/D sky130_fd_sc_hd__or3_1
X_5057_ _4986_/B _5050_/X _5045_/X _5009_/B _5065_/A vssd1 vssd1 vccd1 vccd1 _5064_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_57_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5959_ _5960_/A _5960_/B _5960_/C vssd1 vssd1 vccd1 vccd1 _5961_/A sky130_fd_sc_hd__a21oi_1
XFILLER_25_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8678_ _8681_/CLK _8678_/D vssd1 vssd1 vccd1 vccd1 _8678_/Q sky130_fd_sc_hd__dfxtp_1
X_7629_ _7629_/A vssd1 vssd1 vccd1 vccd1 _7722_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_4_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7980_ _7980_/A _8023_/A _7980_/C vssd1 vssd1 vccd1 vccd1 _8023_/B sky130_fd_sc_hd__nand3_2
XFILLER_54_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6931_ _7336_/S _6931_/B vssd1 vssd1 vccd1 vccd1 _6932_/B sky130_fd_sc_hd__xor2_1
XFILLER_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6862_ _6862_/A _6862_/B vssd1 vssd1 vccd1 vccd1 _6863_/B sky130_fd_sc_hd__and2_1
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8601_ _8671_/CLK _8601_/D vssd1 vssd1 vccd1 vccd1 _8601_/Q sky130_fd_sc_hd__dfxtp_1
X_5813_ _5813_/A _5944_/A vssd1 vssd1 vccd1 vccd1 _5814_/A sky130_fd_sc_hd__and2_1
XFILLER_22_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6793_ _6792_/A _7127_/A _6793_/C vssd1 vssd1 vccd1 vccd1 _6793_/X sky130_fd_sc_hd__and3b_1
X_8532_ _4771_/X _8520_/X _8530_/X _8531_/Y vssd1 vssd1 vccd1 vccd1 _8727_/D sky130_fd_sc_hd__a31oi_1
X_5744_ _5833_/A _6193_/B _5743_/Y vssd1 vssd1 vccd1 vccd1 _5745_/B sky130_fd_sc_hd__o21a_1
X_5675_ _6120_/A _6193_/A _5673_/A _6033_/A vssd1 vssd1 vccd1 vccd1 _6038_/A sky130_fd_sc_hd__o31a_2
X_8463_ _8463_/A _8463_/B vssd1 vssd1 vccd1 vccd1 _8464_/B sky130_fd_sc_hd__xnor2_1
X_7414_ _6880_/X _6892_/B _7414_/S vssd1 vssd1 vccd1 vccd1 _7417_/A sky130_fd_sc_hd__mux2_1
X_4626_ _8594_/Q _4628_/C _4607_/X vssd1 vssd1 vccd1 vccd1 _4626_/Y sky130_fd_sc_hd__o21ai_1
X_8394_ _8394_/A _8394_/B vssd1 vssd1 vccd1 vccd1 _8421_/A sky130_fd_sc_hd__xnor2_1
X_7345_ _7345_/A _7345_/B vssd1 vssd1 vccd1 vccd1 _7382_/A sky130_fd_sc_hd__xnor2_1
X_4557_ _8632_/Q _4563_/B vssd1 vssd1 vccd1 vccd1 _4558_/A sky130_fd_sc_hd__and2_1
XFILLER_103_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7276_ _7275_/A _7276_/B vssd1 vssd1 vccd1 vccd1 _7276_/X sky130_fd_sc_hd__and2b_1
X_4488_ _4848_/A vssd1 vssd1 vccd1 vccd1 _4847_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6227_ _6227_/A _6227_/B vssd1 vssd1 vccd1 vccd1 _6278_/B sky130_fd_sc_hd__nor2_2
XFILLER_97_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6158_ _6303_/A _6094_/A _6303_/B vssd1 vssd1 vccd1 vccd1 _6158_/X sky130_fd_sc_hd__o21a_1
XFILLER_97_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5109_ _5143_/A _5109_/B _5109_/C _5109_/D vssd1 vssd1 vccd1 vccd1 _5109_/X sky130_fd_sc_hd__or4_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6089_ _6089_/A _6089_/B vssd1 vssd1 vccd1 vccd1 _6152_/B sky130_fd_sc_hd__xor2_1
XFILLER_45_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8775__42 vssd1 vssd1 vccd1 vccd1 _8775__42/HI _8870_/A sky130_fd_sc_hd__conb_1
XFILLER_63_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5460_ _5780_/A vssd1 vssd1 vccd1 vccd1 _5872_/A sky130_fd_sc_hd__clkbuf_2
X_4411_ _4413_/A vssd1 vssd1 vccd1 vccd1 _4411_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5391_ _4647_/A _8601_/Q vssd1 vssd1 vccd1 vccd1 _5410_/A sky130_fd_sc_hd__and2b_1
X_7130_ _7130_/A _7130_/B vssd1 vssd1 vccd1 vccd1 _7133_/C sky130_fd_sc_hd__xnor2_1
X_4342_ _4344_/A vssd1 vssd1 vccd1 vccd1 _4342_/Y sky130_fd_sc_hd__inv_2
X_7061_ _7065_/A _7430_/B _6836_/A _7059_/Y _7067_/A vssd1 vssd1 vccd1 vccd1 _7270_/A
+ sky130_fd_sc_hd__o32a_2
XFILLER_98_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6012_ _6161_/B _6012_/B vssd1 vssd1 vccd1 vccd1 _6013_/B sky130_fd_sc_hd__xnor2_1
.ends

