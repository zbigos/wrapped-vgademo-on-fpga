VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_vgademo_on_fpga
  CLASS BLOCK ;
  FOREIGN wrapped_vgademo_on_fpga ;
  ORIGIN 0.000 0.000 ;
  SIZE 300.000 BY 280.000 ;
  PIN active
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.790 276.000 2.350 280.000 ;
    END
  END active
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.150 276.000 9.710 280.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.790 276.000 48.350 280.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.470 276.000 52.030 280.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.610 276.000 56.170 280.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.290 276.000 59.850 280.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.970 276.000 63.530 280.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.110 276.000 67.670 280.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.790 276.000 71.350 280.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.470 276.000 75.030 280.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.610 276.000 79.170 280.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.290 276.000 82.850 280.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.290 276.000 13.850 280.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.970 276.000 86.530 280.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.110 276.000 90.670 280.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.790 276.000 94.350 280.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.470 276.000 98.030 280.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.610 276.000 102.170 280.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.290 276.000 105.850 280.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.430 276.000 109.990 280.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.110 276.000 113.670 280.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.790 276.000 117.350 280.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.930 276.000 121.490 280.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.970 276.000 17.530 280.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.610 276.000 125.170 280.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.290 276.000 128.850 280.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.430 276.000 132.990 280.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.110 276.000 136.670 280.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.790 276.000 140.350 280.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.930 276.000 144.490 280.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.610 276.000 148.170 280.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.750 276.000 152.310 280.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.650 276.000 21.210 280.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.790 276.000 25.350 280.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.470 276.000 29.030 280.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.150 276.000 32.710 280.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.290 276.000 36.850 280.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.970 276.000 40.530 280.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.650 276.000 44.210 280.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 128.940 300.000 130.140 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 169.060 300.000 170.260 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 173.140 300.000 174.340 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 176.540 300.000 177.740 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 180.620 300.000 181.820 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 184.700 300.000 185.900 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 188.780 300.000 189.980 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 192.860 300.000 194.060 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 196.940 300.000 198.140 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 201.020 300.000 202.220 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 205.100 300.000 206.300 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 133.020 300.000 134.220 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 209.180 300.000 210.380 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 212.580 300.000 213.780 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 216.660 300.000 217.860 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 220.740 300.000 221.940 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 224.820 300.000 226.020 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 228.900 300.000 230.100 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 232.980 300.000 234.180 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 237.060 300.000 238.260 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 241.140 300.000 242.340 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 245.220 300.000 246.420 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 137.100 300.000 138.300 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 248.620 300.000 249.820 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 252.700 300.000 253.900 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 256.780 300.000 257.980 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 260.860 300.000 262.060 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 264.940 300.000 266.140 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 269.020 300.000 270.220 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 273.100 300.000 274.300 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 277.180 300.000 278.380 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 141.180 300.000 142.380 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 144.580 300.000 145.780 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 148.660 300.000 149.860 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 152.740 300.000 153.940 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 156.820 300.000 158.020 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 160.900 300.000 162.100 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 164.980 300.000 166.180 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.430 276.000 155.990 280.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.610 276.000 194.170 280.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.750 276.000 198.310 280.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.430 276.000 201.990 280.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.570 276.000 206.130 280.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.250 276.000 209.810 280.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.930 276.000 213.490 280.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.070 276.000 217.630 280.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.750 276.000 221.310 280.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.430 276.000 224.990 280.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.570 276.000 229.130 280.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.110 276.000 159.670 280.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.250 276.000 232.810 280.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.930 276.000 236.490 280.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.070 276.000 240.630 280.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.750 276.000 244.310 280.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.430 276.000 247.990 280.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.570 276.000 252.130 280.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.250 276.000 255.810 280.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.390 276.000 259.950 280.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.070 276.000 263.630 280.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.750 276.000 267.310 280.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.250 276.000 163.810 280.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.890 276.000 271.450 280.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.570 276.000 275.130 280.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.250 276.000 278.810 280.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.390 276.000 282.950 280.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.070 276.000 286.630 280.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.750 276.000 290.310 280.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.890 276.000 294.450 280.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.570 276.000 298.130 280.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.930 276.000 167.490 280.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.610 276.000 171.170 280.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.750 276.000 175.310 280.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.430 276.000 178.990 280.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.110 276.000 182.670 280.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.250 276.000 186.810 280.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.930 276.000 190.490 280.000 ;
    END
  END io_out[9]
  PIN la1_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1.780 4.000 2.980 ;
    END
  END la1_data_in[0]
  PIN la1_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.300 4.000 46.500 ;
    END
  END la1_data_in[10]
  PIN la1_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.380 4.000 50.580 ;
    END
  END la1_data_in[11]
  PIN la1_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.140 4.000 55.340 ;
    END
  END la1_data_in[12]
  PIN la1_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.220 4.000 59.420 ;
    END
  END la1_data_in[13]
  PIN la1_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.980 4.000 64.180 ;
    END
  END la1_data_in[14]
  PIN la1_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 67.060 4.000 68.260 ;
    END
  END la1_data_in[15]
  PIN la1_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.820 4.000 73.020 ;
    END
  END la1_data_in[16]
  PIN la1_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 75.900 4.000 77.100 ;
    END
  END la1_data_in[17]
  PIN la1_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 79.980 4.000 81.180 ;
    END
  END la1_data_in[18]
  PIN la1_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.740 4.000 85.940 ;
    END
  END la1_data_in[19]
  PIN la1_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 5.860 4.000 7.060 ;
    END
  END la1_data_in[1]
  PIN la1_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.820 4.000 90.020 ;
    END
  END la1_data_in[20]
  PIN la1_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.580 4.000 94.780 ;
    END
  END la1_data_in[21]
  PIN la1_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.660 4.000 98.860 ;
    END
  END la1_data_in[22]
  PIN la1_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.420 4.000 103.620 ;
    END
  END la1_data_in[23]
  PIN la1_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.500 4.000 107.700 ;
    END
  END la1_data_in[24]
  PIN la1_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.580 4.000 111.780 ;
    END
  END la1_data_in[25]
  PIN la1_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.340 4.000 116.540 ;
    END
  END la1_data_in[26]
  PIN la1_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.420 4.000 120.620 ;
    END
  END la1_data_in[27]
  PIN la1_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 124.180 4.000 125.380 ;
    END
  END la1_data_in[28]
  PIN la1_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 128.260 4.000 129.460 ;
    END
  END la1_data_in[29]
  PIN la1_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 9.940 4.000 11.140 ;
    END
  END la1_data_in[2]
  PIN la1_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 133.020 4.000 134.220 ;
    END
  END la1_data_in[30]
  PIN la1_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.100 4.000 138.300 ;
    END
  END la1_data_in[31]
  PIN la1_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 14.700 4.000 15.900 ;
    END
  END la1_data_in[3]
  PIN la1_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 18.780 4.000 19.980 ;
    END
  END la1_data_in[4]
  PIN la1_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.540 4.000 24.740 ;
    END
  END la1_data_in[5]
  PIN la1_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.620 4.000 28.820 ;
    END
  END la1_data_in[6]
  PIN la1_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.380 4.000 33.580 ;
    END
  END la1_data_in[7]
  PIN la1_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.460 4.000 37.660 ;
    END
  END la1_data_in[8]
  PIN la1_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.540 4.000 41.740 ;
    END
  END la1_data_in[9]
  PIN la1_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.860 4.000 143.060 ;
    END
  END la1_data_out[0]
  PIN la1_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.380 4.000 186.580 ;
    END
  END la1_data_out[10]
  PIN la1_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.460 4.000 190.660 ;
    END
  END la1_data_out[11]
  PIN la1_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 194.220 4.000 195.420 ;
    END
  END la1_data_out[12]
  PIN la1_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.300 4.000 199.500 ;
    END
  END la1_data_out[13]
  PIN la1_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 203.060 4.000 204.260 ;
    END
  END la1_data_out[14]
  PIN la1_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.140 4.000 208.340 ;
    END
  END la1_data_out[15]
  PIN la1_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 211.900 4.000 213.100 ;
    END
  END la1_data_out[16]
  PIN la1_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 215.980 4.000 217.180 ;
    END
  END la1_data_out[17]
  PIN la1_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 220.060 4.000 221.260 ;
    END
  END la1_data_out[18]
  PIN la1_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.820 4.000 226.020 ;
    END
  END la1_data_out[19]
  PIN la1_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.940 4.000 147.140 ;
    END
  END la1_data_out[1]
  PIN la1_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 228.900 4.000 230.100 ;
    END
  END la1_data_out[20]
  PIN la1_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.660 4.000 234.860 ;
    END
  END la1_data_out[21]
  PIN la1_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 237.740 4.000 238.940 ;
    END
  END la1_data_out[22]
  PIN la1_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.500 4.000 243.700 ;
    END
  END la1_data_out[23]
  PIN la1_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 246.580 4.000 247.780 ;
    END
  END la1_data_out[24]
  PIN la1_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 250.660 4.000 251.860 ;
    END
  END la1_data_out[25]
  PIN la1_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.420 4.000 256.620 ;
    END
  END la1_data_out[26]
  PIN la1_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.500 4.000 260.700 ;
    END
  END la1_data_out[27]
  PIN la1_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 264.260 4.000 265.460 ;
    END
  END la1_data_out[28]
  PIN la1_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 268.340 4.000 269.540 ;
    END
  END la1_data_out[29]
  PIN la1_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 150.020 4.000 151.220 ;
    END
  END la1_data_out[2]
  PIN la1_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 273.100 4.000 274.300 ;
    END
  END la1_data_out[30]
  PIN la1_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 277.180 4.000 278.380 ;
    END
  END la1_data_out[31]
  PIN la1_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 154.780 4.000 155.980 ;
    END
  END la1_data_out[3]
  PIN la1_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 158.860 4.000 160.060 ;
    END
  END la1_data_out[4]
  PIN la1_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.620 4.000 164.820 ;
    END
  END la1_data_out[5]
  PIN la1_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 167.700 4.000 168.900 ;
    END
  END la1_data_out[6]
  PIN la1_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.460 4.000 173.660 ;
    END
  END la1_data_out[7]
  PIN la1_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.540 4.000 177.740 ;
    END
  END la1_data_out[8]
  PIN la1_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.620 4.000 181.820 ;
    END
  END la1_data_out[9]
  PIN la1_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 1.100 300.000 2.300 ;
    END
  END la1_oenb[0]
  PIN la1_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 40.540 300.000 41.740 ;
    END
  END la1_oenb[10]
  PIN la1_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 44.620 300.000 45.820 ;
    END
  END la1_oenb[11]
  PIN la1_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 48.700 300.000 49.900 ;
    END
  END la1_oenb[12]
  PIN la1_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 52.780 300.000 53.980 ;
    END
  END la1_oenb[13]
  PIN la1_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 56.860 300.000 58.060 ;
    END
  END la1_oenb[14]
  PIN la1_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 60.940 300.000 62.140 ;
    END
  END la1_oenb[15]
  PIN la1_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 65.020 300.000 66.220 ;
    END
  END la1_oenb[16]
  PIN la1_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 69.100 300.000 70.300 ;
    END
  END la1_oenb[17]
  PIN la1_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 72.500 300.000 73.700 ;
    END
  END la1_oenb[18]
  PIN la1_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 76.580 300.000 77.780 ;
    END
  END la1_oenb[19]
  PIN la1_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 4.500 300.000 5.700 ;
    END
  END la1_oenb[1]
  PIN la1_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 80.660 300.000 81.860 ;
    END
  END la1_oenb[20]
  PIN la1_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 84.740 300.000 85.940 ;
    END
  END la1_oenb[21]
  PIN la1_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 88.820 300.000 90.020 ;
    END
  END la1_oenb[22]
  PIN la1_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 92.900 300.000 94.100 ;
    END
  END la1_oenb[23]
  PIN la1_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 96.980 300.000 98.180 ;
    END
  END la1_oenb[24]
  PIN la1_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 101.060 300.000 102.260 ;
    END
  END la1_oenb[25]
  PIN la1_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 105.140 300.000 106.340 ;
    END
  END la1_oenb[26]
  PIN la1_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 108.540 300.000 109.740 ;
    END
  END la1_oenb[27]
  PIN la1_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 112.620 300.000 113.820 ;
    END
  END la1_oenb[28]
  PIN la1_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 116.700 300.000 117.900 ;
    END
  END la1_oenb[29]
  PIN la1_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 8.580 300.000 9.780 ;
    END
  END la1_oenb[2]
  PIN la1_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 120.780 300.000 121.980 ;
    END
  END la1_oenb[30]
  PIN la1_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 124.860 300.000 126.060 ;
    END
  END la1_oenb[31]
  PIN la1_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 12.660 300.000 13.860 ;
    END
  END la1_oenb[3]
  PIN la1_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 16.740 300.000 17.940 ;
    END
  END la1_oenb[4]
  PIN la1_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 20.820 300.000 22.020 ;
    END
  END la1_oenb[5]
  PIN la1_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 24.900 300.000 26.100 ;
    END
  END la1_oenb[6]
  PIN la1_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 28.980 300.000 30.180 ;
    END
  END la1_oenb[7]
  PIN la1_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 33.060 300.000 34.260 ;
    END
  END la1_oenb[8]
  PIN la1_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 36.460 300.000 37.660 ;
    END
  END la1_oenb[9]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 2.480 22.640 266.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 2.480 176.240 266.800 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 2.480 99.440 266.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 2.480 253.040 266.800 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.470 276.000 6.030 280.000 ;
    END
  END wb_clk_i
  OBS
      LAYER li1 ;
        RECT 5.520 2.635 294.400 266.645 ;
      LAYER met1 ;
        RECT 1.910 2.480 298.010 271.960 ;
      LAYER met2 ;
        RECT 2.630 275.720 5.190 277.965 ;
        RECT 6.310 275.720 8.870 277.965 ;
        RECT 9.990 275.720 13.010 277.965 ;
        RECT 14.130 275.720 16.690 277.965 ;
        RECT 17.810 275.720 20.370 277.965 ;
        RECT 21.490 275.720 24.510 277.965 ;
        RECT 25.630 275.720 28.190 277.965 ;
        RECT 29.310 275.720 31.870 277.965 ;
        RECT 32.990 275.720 36.010 277.965 ;
        RECT 37.130 275.720 39.690 277.965 ;
        RECT 40.810 275.720 43.370 277.965 ;
        RECT 44.490 275.720 47.510 277.965 ;
        RECT 48.630 275.720 51.190 277.965 ;
        RECT 52.310 275.720 55.330 277.965 ;
        RECT 56.450 275.720 59.010 277.965 ;
        RECT 60.130 275.720 62.690 277.965 ;
        RECT 63.810 275.720 66.830 277.965 ;
        RECT 67.950 275.720 70.510 277.965 ;
        RECT 71.630 275.720 74.190 277.965 ;
        RECT 75.310 275.720 78.330 277.965 ;
        RECT 79.450 275.720 82.010 277.965 ;
        RECT 83.130 275.720 85.690 277.965 ;
        RECT 86.810 275.720 89.830 277.965 ;
        RECT 90.950 275.720 93.510 277.965 ;
        RECT 94.630 275.720 97.190 277.965 ;
        RECT 98.310 275.720 101.330 277.965 ;
        RECT 102.450 275.720 105.010 277.965 ;
        RECT 106.130 275.720 109.150 277.965 ;
        RECT 110.270 275.720 112.830 277.965 ;
        RECT 113.950 275.720 116.510 277.965 ;
        RECT 117.630 275.720 120.650 277.965 ;
        RECT 121.770 275.720 124.330 277.965 ;
        RECT 125.450 275.720 128.010 277.965 ;
        RECT 129.130 275.720 132.150 277.965 ;
        RECT 133.270 275.720 135.830 277.965 ;
        RECT 136.950 275.720 139.510 277.965 ;
        RECT 140.630 275.720 143.650 277.965 ;
        RECT 144.770 275.720 147.330 277.965 ;
        RECT 148.450 275.720 151.470 277.965 ;
        RECT 152.590 275.720 155.150 277.965 ;
        RECT 156.270 275.720 158.830 277.965 ;
        RECT 159.950 275.720 162.970 277.965 ;
        RECT 164.090 275.720 166.650 277.965 ;
        RECT 167.770 275.720 170.330 277.965 ;
        RECT 171.450 275.720 174.470 277.965 ;
        RECT 175.590 275.720 178.150 277.965 ;
        RECT 179.270 275.720 181.830 277.965 ;
        RECT 182.950 275.720 185.970 277.965 ;
        RECT 187.090 275.720 189.650 277.965 ;
        RECT 190.770 275.720 193.330 277.965 ;
        RECT 194.450 275.720 197.470 277.965 ;
        RECT 198.590 275.720 201.150 277.965 ;
        RECT 202.270 275.720 205.290 277.965 ;
        RECT 206.410 275.720 208.970 277.965 ;
        RECT 210.090 275.720 212.650 277.965 ;
        RECT 213.770 275.720 216.790 277.965 ;
        RECT 217.910 275.720 220.470 277.965 ;
        RECT 221.590 275.720 224.150 277.965 ;
        RECT 225.270 275.720 228.290 277.965 ;
        RECT 229.410 275.720 231.970 277.965 ;
        RECT 233.090 275.720 235.650 277.965 ;
        RECT 236.770 275.720 239.790 277.965 ;
        RECT 240.910 275.720 243.470 277.965 ;
        RECT 244.590 275.720 247.150 277.965 ;
        RECT 248.270 275.720 251.290 277.965 ;
        RECT 252.410 275.720 254.970 277.965 ;
        RECT 256.090 275.720 259.110 277.965 ;
        RECT 260.230 275.720 262.790 277.965 ;
        RECT 263.910 275.720 266.470 277.965 ;
        RECT 267.590 275.720 270.610 277.965 ;
        RECT 271.730 275.720 274.290 277.965 ;
        RECT 275.410 275.720 277.970 277.965 ;
        RECT 279.090 275.720 282.110 277.965 ;
        RECT 283.230 275.720 285.790 277.965 ;
        RECT 286.910 275.720 289.470 277.965 ;
        RECT 290.590 275.720 293.610 277.965 ;
        RECT 294.730 275.720 297.290 277.965 ;
        RECT 1.940 2.480 297.980 275.720 ;
      LAYER met3 ;
        RECT 4.400 276.780 295.600 277.945 ;
        RECT 4.000 274.700 296.000 276.780 ;
        RECT 4.400 272.700 295.600 274.700 ;
        RECT 4.000 270.620 296.000 272.700 ;
        RECT 4.000 269.940 295.600 270.620 ;
        RECT 4.400 268.620 295.600 269.940 ;
        RECT 4.400 267.940 296.000 268.620 ;
        RECT 4.000 266.540 296.000 267.940 ;
        RECT 4.000 265.860 295.600 266.540 ;
        RECT 4.400 264.540 295.600 265.860 ;
        RECT 4.400 263.860 296.000 264.540 ;
        RECT 4.000 262.460 296.000 263.860 ;
        RECT 4.000 261.100 295.600 262.460 ;
        RECT 4.400 260.460 295.600 261.100 ;
        RECT 4.400 259.100 296.000 260.460 ;
        RECT 4.000 258.380 296.000 259.100 ;
        RECT 4.000 257.020 295.600 258.380 ;
        RECT 4.400 256.380 295.600 257.020 ;
        RECT 4.400 255.020 296.000 256.380 ;
        RECT 4.000 254.300 296.000 255.020 ;
        RECT 4.000 252.300 295.600 254.300 ;
        RECT 4.000 252.260 296.000 252.300 ;
        RECT 4.400 250.260 296.000 252.260 ;
        RECT 4.000 250.220 296.000 250.260 ;
        RECT 4.000 248.220 295.600 250.220 ;
        RECT 4.000 248.180 296.000 248.220 ;
        RECT 4.400 246.820 296.000 248.180 ;
        RECT 4.400 246.180 295.600 246.820 ;
        RECT 4.000 244.820 295.600 246.180 ;
        RECT 4.000 244.100 296.000 244.820 ;
        RECT 4.400 242.740 296.000 244.100 ;
        RECT 4.400 242.100 295.600 242.740 ;
        RECT 4.000 240.740 295.600 242.100 ;
        RECT 4.000 239.340 296.000 240.740 ;
        RECT 4.400 238.660 296.000 239.340 ;
        RECT 4.400 237.340 295.600 238.660 ;
        RECT 4.000 236.660 295.600 237.340 ;
        RECT 4.000 235.260 296.000 236.660 ;
        RECT 4.400 234.580 296.000 235.260 ;
        RECT 4.400 233.260 295.600 234.580 ;
        RECT 4.000 232.580 295.600 233.260 ;
        RECT 4.000 230.500 296.000 232.580 ;
        RECT 4.400 228.500 295.600 230.500 ;
        RECT 4.000 226.420 296.000 228.500 ;
        RECT 4.400 224.420 295.600 226.420 ;
        RECT 4.000 222.340 296.000 224.420 ;
        RECT 4.000 221.660 295.600 222.340 ;
        RECT 4.400 220.340 295.600 221.660 ;
        RECT 4.400 219.660 296.000 220.340 ;
        RECT 4.000 218.260 296.000 219.660 ;
        RECT 4.000 217.580 295.600 218.260 ;
        RECT 4.400 216.260 295.600 217.580 ;
        RECT 4.400 215.580 296.000 216.260 ;
        RECT 4.000 214.180 296.000 215.580 ;
        RECT 4.000 213.500 295.600 214.180 ;
        RECT 4.400 212.180 295.600 213.500 ;
        RECT 4.400 211.500 296.000 212.180 ;
        RECT 4.000 210.780 296.000 211.500 ;
        RECT 4.000 208.780 295.600 210.780 ;
        RECT 4.000 208.740 296.000 208.780 ;
        RECT 4.400 206.740 296.000 208.740 ;
        RECT 4.000 206.700 296.000 206.740 ;
        RECT 4.000 204.700 295.600 206.700 ;
        RECT 4.000 204.660 296.000 204.700 ;
        RECT 4.400 202.660 296.000 204.660 ;
        RECT 4.000 202.620 296.000 202.660 ;
        RECT 4.000 200.620 295.600 202.620 ;
        RECT 4.000 199.900 296.000 200.620 ;
        RECT 4.400 198.540 296.000 199.900 ;
        RECT 4.400 197.900 295.600 198.540 ;
        RECT 4.000 196.540 295.600 197.900 ;
        RECT 4.000 195.820 296.000 196.540 ;
        RECT 4.400 194.460 296.000 195.820 ;
        RECT 4.400 193.820 295.600 194.460 ;
        RECT 4.000 192.460 295.600 193.820 ;
        RECT 4.000 191.060 296.000 192.460 ;
        RECT 4.400 190.380 296.000 191.060 ;
        RECT 4.400 189.060 295.600 190.380 ;
        RECT 4.000 188.380 295.600 189.060 ;
        RECT 4.000 186.980 296.000 188.380 ;
        RECT 4.400 186.300 296.000 186.980 ;
        RECT 4.400 184.980 295.600 186.300 ;
        RECT 4.000 184.300 295.600 184.980 ;
        RECT 4.000 182.220 296.000 184.300 ;
        RECT 4.400 180.220 295.600 182.220 ;
        RECT 4.000 178.140 296.000 180.220 ;
        RECT 4.400 176.140 295.600 178.140 ;
        RECT 4.000 174.740 296.000 176.140 ;
        RECT 4.000 174.060 295.600 174.740 ;
        RECT 4.400 172.740 295.600 174.060 ;
        RECT 4.400 172.060 296.000 172.740 ;
        RECT 4.000 170.660 296.000 172.060 ;
        RECT 4.000 169.300 295.600 170.660 ;
        RECT 4.400 168.660 295.600 169.300 ;
        RECT 4.400 167.300 296.000 168.660 ;
        RECT 4.000 166.580 296.000 167.300 ;
        RECT 4.000 165.220 295.600 166.580 ;
        RECT 4.400 164.580 295.600 165.220 ;
        RECT 4.400 163.220 296.000 164.580 ;
        RECT 4.000 162.500 296.000 163.220 ;
        RECT 4.000 160.500 295.600 162.500 ;
        RECT 4.000 160.460 296.000 160.500 ;
        RECT 4.400 158.460 296.000 160.460 ;
        RECT 4.000 158.420 296.000 158.460 ;
        RECT 4.000 156.420 295.600 158.420 ;
        RECT 4.000 156.380 296.000 156.420 ;
        RECT 4.400 154.380 296.000 156.380 ;
        RECT 4.000 154.340 296.000 154.380 ;
        RECT 4.000 152.340 295.600 154.340 ;
        RECT 4.000 151.620 296.000 152.340 ;
        RECT 4.400 150.260 296.000 151.620 ;
        RECT 4.400 149.620 295.600 150.260 ;
        RECT 4.000 148.260 295.600 149.620 ;
        RECT 4.000 147.540 296.000 148.260 ;
        RECT 4.400 146.180 296.000 147.540 ;
        RECT 4.400 145.540 295.600 146.180 ;
        RECT 4.000 144.180 295.600 145.540 ;
        RECT 4.000 143.460 296.000 144.180 ;
        RECT 4.400 142.780 296.000 143.460 ;
        RECT 4.400 141.460 295.600 142.780 ;
        RECT 4.000 140.780 295.600 141.460 ;
        RECT 4.000 138.700 296.000 140.780 ;
        RECT 4.400 136.700 295.600 138.700 ;
        RECT 4.000 134.620 296.000 136.700 ;
        RECT 4.400 132.620 295.600 134.620 ;
        RECT 4.000 130.540 296.000 132.620 ;
        RECT 4.000 129.860 295.600 130.540 ;
        RECT 4.400 128.540 295.600 129.860 ;
        RECT 4.400 127.860 296.000 128.540 ;
        RECT 4.000 126.460 296.000 127.860 ;
        RECT 4.000 125.780 295.600 126.460 ;
        RECT 4.400 124.460 295.600 125.780 ;
        RECT 4.400 123.780 296.000 124.460 ;
        RECT 4.000 122.380 296.000 123.780 ;
        RECT 4.000 121.020 295.600 122.380 ;
        RECT 4.400 120.380 295.600 121.020 ;
        RECT 4.400 119.020 296.000 120.380 ;
        RECT 4.000 118.300 296.000 119.020 ;
        RECT 4.000 116.940 295.600 118.300 ;
        RECT 4.400 116.300 295.600 116.940 ;
        RECT 4.400 114.940 296.000 116.300 ;
        RECT 4.000 114.220 296.000 114.940 ;
        RECT 4.000 112.220 295.600 114.220 ;
        RECT 4.000 112.180 296.000 112.220 ;
        RECT 4.400 110.180 296.000 112.180 ;
        RECT 4.000 110.140 296.000 110.180 ;
        RECT 4.000 108.140 295.600 110.140 ;
        RECT 4.000 108.100 296.000 108.140 ;
        RECT 4.400 106.740 296.000 108.100 ;
        RECT 4.400 106.100 295.600 106.740 ;
        RECT 4.000 104.740 295.600 106.100 ;
        RECT 4.000 104.020 296.000 104.740 ;
        RECT 4.400 102.660 296.000 104.020 ;
        RECT 4.400 102.020 295.600 102.660 ;
        RECT 4.000 100.660 295.600 102.020 ;
        RECT 4.000 99.260 296.000 100.660 ;
        RECT 4.400 98.580 296.000 99.260 ;
        RECT 4.400 97.260 295.600 98.580 ;
        RECT 4.000 96.580 295.600 97.260 ;
        RECT 4.000 95.180 296.000 96.580 ;
        RECT 4.400 94.500 296.000 95.180 ;
        RECT 4.400 93.180 295.600 94.500 ;
        RECT 4.000 92.500 295.600 93.180 ;
        RECT 4.000 90.420 296.000 92.500 ;
        RECT 4.400 88.420 295.600 90.420 ;
        RECT 4.000 86.340 296.000 88.420 ;
        RECT 4.400 84.340 295.600 86.340 ;
        RECT 4.000 82.260 296.000 84.340 ;
        RECT 4.000 81.580 295.600 82.260 ;
        RECT 4.400 80.260 295.600 81.580 ;
        RECT 4.400 79.580 296.000 80.260 ;
        RECT 4.000 78.180 296.000 79.580 ;
        RECT 4.000 77.500 295.600 78.180 ;
        RECT 4.400 76.180 295.600 77.500 ;
        RECT 4.400 75.500 296.000 76.180 ;
        RECT 4.000 74.100 296.000 75.500 ;
        RECT 4.000 73.420 295.600 74.100 ;
        RECT 4.400 72.100 295.600 73.420 ;
        RECT 4.400 71.420 296.000 72.100 ;
        RECT 4.000 70.700 296.000 71.420 ;
        RECT 4.000 68.700 295.600 70.700 ;
        RECT 4.000 68.660 296.000 68.700 ;
        RECT 4.400 66.660 296.000 68.660 ;
        RECT 4.000 66.620 296.000 66.660 ;
        RECT 4.000 64.620 295.600 66.620 ;
        RECT 4.000 64.580 296.000 64.620 ;
        RECT 4.400 62.580 296.000 64.580 ;
        RECT 4.000 62.540 296.000 62.580 ;
        RECT 4.000 60.540 295.600 62.540 ;
        RECT 4.000 59.820 296.000 60.540 ;
        RECT 4.400 58.460 296.000 59.820 ;
        RECT 4.400 57.820 295.600 58.460 ;
        RECT 4.000 56.460 295.600 57.820 ;
        RECT 4.000 55.740 296.000 56.460 ;
        RECT 4.400 54.380 296.000 55.740 ;
        RECT 4.400 53.740 295.600 54.380 ;
        RECT 4.000 52.380 295.600 53.740 ;
        RECT 4.000 50.980 296.000 52.380 ;
        RECT 4.400 50.300 296.000 50.980 ;
        RECT 4.400 48.980 295.600 50.300 ;
        RECT 4.000 48.300 295.600 48.980 ;
        RECT 4.000 46.900 296.000 48.300 ;
        RECT 4.400 46.220 296.000 46.900 ;
        RECT 4.400 44.900 295.600 46.220 ;
        RECT 4.000 44.220 295.600 44.900 ;
        RECT 4.000 42.140 296.000 44.220 ;
        RECT 4.400 40.140 295.600 42.140 ;
        RECT 4.000 38.060 296.000 40.140 ;
        RECT 4.400 36.060 295.600 38.060 ;
        RECT 4.000 34.660 296.000 36.060 ;
        RECT 4.000 33.980 295.600 34.660 ;
        RECT 4.400 32.660 295.600 33.980 ;
        RECT 4.400 31.980 296.000 32.660 ;
        RECT 4.000 30.580 296.000 31.980 ;
        RECT 4.000 29.220 295.600 30.580 ;
        RECT 4.400 28.580 295.600 29.220 ;
        RECT 4.400 27.220 296.000 28.580 ;
        RECT 4.000 26.500 296.000 27.220 ;
        RECT 4.000 25.140 295.600 26.500 ;
        RECT 4.400 24.500 295.600 25.140 ;
        RECT 4.400 23.140 296.000 24.500 ;
        RECT 4.000 22.420 296.000 23.140 ;
        RECT 4.000 20.420 295.600 22.420 ;
        RECT 4.000 20.380 296.000 20.420 ;
        RECT 4.400 18.380 296.000 20.380 ;
        RECT 4.000 18.340 296.000 18.380 ;
        RECT 4.000 16.340 295.600 18.340 ;
        RECT 4.000 16.300 296.000 16.340 ;
        RECT 4.400 14.300 296.000 16.300 ;
        RECT 4.000 14.260 296.000 14.300 ;
        RECT 4.000 12.260 295.600 14.260 ;
        RECT 4.000 11.540 296.000 12.260 ;
        RECT 4.400 10.180 296.000 11.540 ;
        RECT 4.400 9.540 295.600 10.180 ;
        RECT 4.000 8.180 295.600 9.540 ;
        RECT 4.000 7.460 296.000 8.180 ;
        RECT 4.400 6.100 296.000 7.460 ;
        RECT 4.400 5.460 295.600 6.100 ;
        RECT 4.000 4.100 295.600 5.460 ;
        RECT 4.000 3.380 296.000 4.100 ;
        RECT 4.400 2.700 296.000 3.380 ;
        RECT 4.400 2.555 295.600 2.700 ;
      LAYER met4 ;
        RECT 7.655 267.200 281.225 271.145 ;
        RECT 7.655 71.575 20.640 267.200 ;
        RECT 23.040 71.575 97.440 267.200 ;
        RECT 99.840 71.575 174.240 267.200 ;
        RECT 176.640 71.575 251.040 267.200 ;
        RECT 253.440 71.575 281.225 267.200 ;
  END
END wrapped_vgademo_on_fpga
END LIBRARY

