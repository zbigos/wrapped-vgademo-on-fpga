VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_vgademo_on_fpga
  CLASS BLOCK ;
  FOREIGN wrapped_vgademo_on_fpga ;
  ORIGIN 0.000 0.000 ;
  SIZE 300.000 BY 300.000 ;
  PIN active
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.710 296.000 3.270 300.000 ;
    END
  END active
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.210 296.000 14.770 300.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.090 296.000 73.650 300.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.070 296.000 79.630 300.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.590 296.000 85.150 300.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.570 296.000 91.130 300.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.550 296.000 97.110 300.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.530 296.000 103.090 300.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.510 296.000 109.070 300.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.030 296.000 114.590 300.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.010 296.000 120.570 300.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.990 296.000 126.550 300.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.190 296.000 20.750 300.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.970 296.000 132.530 300.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.950 296.000 138.510 300.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.470 296.000 144.030 300.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.450 296.000 150.010 300.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.430 296.000 155.990 300.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.410 296.000 161.970 300.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.930 296.000 167.490 300.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.910 296.000 173.470 300.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.890 296.000 179.450 300.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.870 296.000 185.430 300.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.170 296.000 26.730 300.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.850 296.000 191.410 300.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.370 296.000 196.930 300.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.350 296.000 202.910 300.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.330 296.000 208.890 300.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.310 296.000 214.870 300.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.290 296.000 220.850 300.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.810 296.000 226.370 300.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.790 296.000 232.350 300.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.690 296.000 32.250 300.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.670 296.000 38.230 300.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.650 296.000 44.210 300.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.630 296.000 50.190 300.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.610 296.000 56.170 300.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.130 296.000 61.690 300.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.110 296.000 67.670 300.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 122.140 300.000 123.340 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 160.220 300.000 161.420 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 164.300 300.000 165.500 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 167.700 300.000 168.900 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 171.780 300.000 172.980 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 175.180 300.000 176.380 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 179.260 300.000 180.460 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 182.660 300.000 183.860 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 186.740 300.000 187.940 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 190.820 300.000 192.020 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 194.220 300.000 195.420 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 126.220 300.000 127.420 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 198.300 300.000 199.500 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 201.700 300.000 202.900 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 205.780 300.000 206.980 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 209.860 300.000 211.060 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 213.260 300.000 214.460 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 217.340 300.000 218.540 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 220.740 300.000 221.940 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 224.820 300.000 226.020 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 228.220 300.000 229.420 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 232.300 300.000 233.500 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 129.620 300.000 130.820 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 236.380 300.000 237.580 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 239.780 300.000 240.980 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 243.860 300.000 245.060 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 247.260 300.000 248.460 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 251.340 300.000 252.540 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 255.420 300.000 256.620 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 258.820 300.000 260.020 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 262.900 300.000 264.100 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 133.700 300.000 134.900 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 137.100 300.000 138.300 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 141.180 300.000 142.380 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 145.260 300.000 146.460 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 148.660 300.000 149.860 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 152.740 300.000 153.940 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 156.140 300.000 157.340 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 266.300 300.000 267.500 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 268.340 4.000 269.540 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 277.860 300.000 279.060 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 281.940 300.000 283.140 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 285.340 300.000 286.540 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.890 0.000 64.450 4.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.250 296.000 255.810 300.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.420 4.000 273.620 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 289.420 300.000 290.620 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.230 296.000 261.790 300.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.210 296.000 267.770 300.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 270.380 300.000 271.580 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.190 296.000 273.750 300.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.670 0.000 107.230 4.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 276.500 4.000 277.700 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.450 0.000 150.010 4.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.710 296.000 279.270 300.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 292.820 300.000 294.020 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 280.580 4.000 281.780 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.230 0.000 192.790 4.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.010 0.000 235.570 4.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 296.900 300.000 298.100 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 256.780 4.000 257.980 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.690 296.000 285.250 300.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.670 296.000 291.230 300.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.660 4.000 285.860 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 288.740 4.000 289.940 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.820 4.000 294.020 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.650 296.000 297.210 300.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 296.900 4.000 298.100 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.790 0.000 278.350 4.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 260.860 4.000 262.060 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.770 296.000 238.330 300.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 264.940 4.000 266.140 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.750 296.000 244.310 300.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.270 296.000 249.830 300.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.110 0.000 21.670 4.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 273.780 300.000 274.980 ;
    END
  END io_out[9]
  PIN la1_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1.100 4.000 2.300 ;
    END
  END la1_data_in[0]
  PIN la1_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.540 4.000 41.740 ;
    END
  END la1_data_in[10]
  PIN la1_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.620 4.000 45.820 ;
    END
  END la1_data_in[11]
  PIN la1_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.700 4.000 49.900 ;
    END
  END la1_data_in[12]
  PIN la1_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 52.780 4.000 53.980 ;
    END
  END la1_data_in[13]
  PIN la1_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 56.860 4.000 58.060 ;
    END
  END la1_data_in[14]
  PIN la1_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 60.940 4.000 62.140 ;
    END
  END la1_data_in[15]
  PIN la1_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.020 4.000 66.220 ;
    END
  END la1_data_in[16]
  PIN la1_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.420 4.000 69.620 ;
    END
  END la1_data_in[17]
  PIN la1_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.500 4.000 73.700 ;
    END
  END la1_data_in[18]
  PIN la1_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.580 4.000 77.780 ;
    END
  END la1_data_in[19]
  PIN la1_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.500 4.000 5.700 ;
    END
  END la1_data_in[1]
  PIN la1_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.660 4.000 81.860 ;
    END
  END la1_data_in[20]
  PIN la1_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.740 4.000 85.940 ;
    END
  END la1_data_in[21]
  PIN la1_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.820 4.000 90.020 ;
    END
  END la1_data_in[22]
  PIN la1_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.900 4.000 94.100 ;
    END
  END la1_data_in[23]
  PIN la1_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.980 4.000 98.180 ;
    END
  END la1_data_in[24]
  PIN la1_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 101.060 4.000 102.260 ;
    END
  END la1_data_in[25]
  PIN la1_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.460 4.000 105.660 ;
    END
  END la1_data_in[26]
  PIN la1_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.540 4.000 109.740 ;
    END
  END la1_data_in[27]
  PIN la1_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.620 4.000 113.820 ;
    END
  END la1_data_in[28]
  PIN la1_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 116.700 4.000 117.900 ;
    END
  END la1_data_in[29]
  PIN la1_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.580 4.000 9.780 ;
    END
  END la1_data_in[2]
  PIN la1_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 120.780 4.000 121.980 ;
    END
  END la1_data_in[30]
  PIN la1_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 124.860 4.000 126.060 ;
    END
  END la1_data_in[31]
  PIN la1_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.660 4.000 13.860 ;
    END
  END la1_data_in[3]
  PIN la1_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.740 4.000 17.940 ;
    END
  END la1_data_in[4]
  PIN la1_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.820 4.000 22.020 ;
    END
  END la1_data_in[5]
  PIN la1_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.900 4.000 26.100 ;
    END
  END la1_data_in[6]
  PIN la1_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.980 4.000 30.180 ;
    END
  END la1_data_in[7]
  PIN la1_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.060 4.000 34.260 ;
    END
  END la1_data_in[8]
  PIN la1_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.460 4.000 37.660 ;
    END
  END la1_data_in[9]
  PIN la1_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 128.940 4.000 130.140 ;
    END
  END la1_data_out[0]
  PIN la1_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.380 4.000 169.580 ;
    END
  END la1_data_out[10]
  PIN la1_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.460 4.000 173.660 ;
    END
  END la1_data_out[11]
  PIN la1_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.540 4.000 177.740 ;
    END
  END la1_data_out[12]
  PIN la1_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.620 4.000 181.820 ;
    END
  END la1_data_out[13]
  PIN la1_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 184.700 4.000 185.900 ;
    END
  END la1_data_out[14]
  PIN la1_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 188.780 4.000 189.980 ;
    END
  END la1_data_out[15]
  PIN la1_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 192.860 4.000 194.060 ;
    END
  END la1_data_out[16]
  PIN la1_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 196.940 4.000 198.140 ;
    END
  END la1_data_out[17]
  PIN la1_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 201.020 4.000 202.220 ;
    END
  END la1_data_out[18]
  PIN la1_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.420 4.000 205.620 ;
    END
  END la1_data_out[19]
  PIN la1_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 133.020 4.000 134.220 ;
    END
  END la1_data_out[1]
  PIN la1_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.500 4.000 209.700 ;
    END
  END la1_data_out[20]
  PIN la1_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.580 4.000 213.780 ;
    END
  END la1_data_out[21]
  PIN la1_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.660 4.000 217.860 ;
    END
  END la1_data_out[22]
  PIN la1_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 220.740 4.000 221.940 ;
    END
  END la1_data_out[23]
  PIN la1_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.820 4.000 226.020 ;
    END
  END la1_data_out[24]
  PIN la1_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 228.900 4.000 230.100 ;
    END
  END la1_data_out[25]
  PIN la1_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 232.980 4.000 234.180 ;
    END
  END la1_data_out[26]
  PIN la1_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.380 4.000 237.580 ;
    END
  END la1_data_out[27]
  PIN la1_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.460 4.000 241.660 ;
    END
  END la1_data_out[28]
  PIN la1_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.540 4.000 245.740 ;
    END
  END la1_data_out[29]
  PIN la1_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.420 4.000 137.620 ;
    END
  END la1_data_out[2]
  PIN la1_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.620 4.000 249.820 ;
    END
  END la1_data_out[30]
  PIN la1_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 252.700 4.000 253.900 ;
    END
  END la1_data_out[31]
  PIN la1_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.500 4.000 141.700 ;
    END
  END la1_data_out[3]
  PIN la1_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.580 4.000 145.780 ;
    END
  END la1_data_out[4]
  PIN la1_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.660 4.000 149.860 ;
    END
  END la1_data_out[5]
  PIN la1_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.740 4.000 153.940 ;
    END
  END la1_data_out[6]
  PIN la1_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.820 4.000 158.020 ;
    END
  END la1_data_out[7]
  PIN la1_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.900 4.000 162.100 ;
    END
  END la1_data_out[8]
  PIN la1_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.980 4.000 166.180 ;
    END
  END la1_data_out[9]
  PIN la1_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 1.100 300.000 2.300 ;
    END
  END la1_oenb[0]
  PIN la1_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 38.500 300.000 39.700 ;
    END
  END la1_oenb[10]
  PIN la1_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 42.580 300.000 43.780 ;
    END
  END la1_oenb[11]
  PIN la1_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 45.980 300.000 47.180 ;
    END
  END la1_oenb[12]
  PIN la1_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 50.060 300.000 51.260 ;
    END
  END la1_oenb[13]
  PIN la1_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 54.140 300.000 55.340 ;
    END
  END la1_oenb[14]
  PIN la1_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 57.540 300.000 58.740 ;
    END
  END la1_oenb[15]
  PIN la1_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 61.620 300.000 62.820 ;
    END
  END la1_oenb[16]
  PIN la1_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 65.020 300.000 66.220 ;
    END
  END la1_oenb[17]
  PIN la1_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 69.100 300.000 70.300 ;
    END
  END la1_oenb[18]
  PIN la1_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 73.180 300.000 74.380 ;
    END
  END la1_oenb[19]
  PIN la1_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 4.500 300.000 5.700 ;
    END
  END la1_oenb[1]
  PIN la1_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 76.580 300.000 77.780 ;
    END
  END la1_oenb[20]
  PIN la1_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 80.660 300.000 81.860 ;
    END
  END la1_oenb[21]
  PIN la1_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 84.060 300.000 85.260 ;
    END
  END la1_oenb[22]
  PIN la1_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 88.140 300.000 89.340 ;
    END
  END la1_oenb[23]
  PIN la1_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 91.540 300.000 92.740 ;
    END
  END la1_oenb[24]
  PIN la1_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 95.620 300.000 96.820 ;
    END
  END la1_oenb[25]
  PIN la1_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 99.700 300.000 100.900 ;
    END
  END la1_oenb[26]
  PIN la1_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 103.100 300.000 104.300 ;
    END
  END la1_oenb[27]
  PIN la1_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 107.180 300.000 108.380 ;
    END
  END la1_oenb[28]
  PIN la1_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 110.580 300.000 111.780 ;
    END
  END la1_oenb[29]
  PIN la1_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 8.580 300.000 9.780 ;
    END
  END la1_oenb[2]
  PIN la1_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 114.660 300.000 115.860 ;
    END
  END la1_oenb[30]
  PIN la1_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 118.740 300.000 119.940 ;
    END
  END la1_oenb[31]
  PIN la1_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 11.980 300.000 13.180 ;
    END
  END la1_oenb[3]
  PIN la1_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 16.060 300.000 17.260 ;
    END
  END la1_oenb[4]
  PIN la1_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 19.460 300.000 20.660 ;
    END
  END la1_oenb[5]
  PIN la1_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 23.540 300.000 24.740 ;
    END
  END la1_oenb[6]
  PIN la1_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 27.620 300.000 28.820 ;
    END
  END la1_oenb[7]
  PIN la1_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 31.020 300.000 32.220 ;
    END
  END la1_oenb[8]
  PIN la1_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 35.100 300.000 36.300 ;
    END
  END la1_oenb[9]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 2.480 22.640 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 2.480 176.240 288.560 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 2.480 99.440 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 2.480 253.040 288.560 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.230 296.000 8.790 300.000 ;
    END
  END wb_clk_i
  OBS
      LAYER li1 ;
        RECT 5.520 2.635 294.400 288.405 ;
      LAYER met1 ;
        RECT 2.830 2.080 297.090 289.640 ;
      LAYER met2 ;
        RECT 3.550 295.720 7.950 297.685 ;
        RECT 9.070 295.720 13.930 297.685 ;
        RECT 15.050 295.720 19.910 297.685 ;
        RECT 21.030 295.720 25.890 297.685 ;
        RECT 27.010 295.720 31.410 297.685 ;
        RECT 32.530 295.720 37.390 297.685 ;
        RECT 38.510 295.720 43.370 297.685 ;
        RECT 44.490 295.720 49.350 297.685 ;
        RECT 50.470 295.720 55.330 297.685 ;
        RECT 56.450 295.720 60.850 297.685 ;
        RECT 61.970 295.720 66.830 297.685 ;
        RECT 67.950 295.720 72.810 297.685 ;
        RECT 73.930 295.720 78.790 297.685 ;
        RECT 79.910 295.720 84.310 297.685 ;
        RECT 85.430 295.720 90.290 297.685 ;
        RECT 91.410 295.720 96.270 297.685 ;
        RECT 97.390 295.720 102.250 297.685 ;
        RECT 103.370 295.720 108.230 297.685 ;
        RECT 109.350 295.720 113.750 297.685 ;
        RECT 114.870 295.720 119.730 297.685 ;
        RECT 120.850 295.720 125.710 297.685 ;
        RECT 126.830 295.720 131.690 297.685 ;
        RECT 132.810 295.720 137.670 297.685 ;
        RECT 138.790 295.720 143.190 297.685 ;
        RECT 144.310 295.720 149.170 297.685 ;
        RECT 150.290 295.720 155.150 297.685 ;
        RECT 156.270 295.720 161.130 297.685 ;
        RECT 162.250 295.720 166.650 297.685 ;
        RECT 167.770 295.720 172.630 297.685 ;
        RECT 173.750 295.720 178.610 297.685 ;
        RECT 179.730 295.720 184.590 297.685 ;
        RECT 185.710 295.720 190.570 297.685 ;
        RECT 191.690 295.720 196.090 297.685 ;
        RECT 197.210 295.720 202.070 297.685 ;
        RECT 203.190 295.720 208.050 297.685 ;
        RECT 209.170 295.720 214.030 297.685 ;
        RECT 215.150 295.720 220.010 297.685 ;
        RECT 221.130 295.720 225.530 297.685 ;
        RECT 226.650 295.720 231.510 297.685 ;
        RECT 232.630 295.720 237.490 297.685 ;
        RECT 238.610 295.720 243.470 297.685 ;
        RECT 244.590 295.720 248.990 297.685 ;
        RECT 250.110 295.720 254.970 297.685 ;
        RECT 256.090 295.720 260.950 297.685 ;
        RECT 262.070 295.720 266.930 297.685 ;
        RECT 268.050 295.720 272.910 297.685 ;
        RECT 274.030 295.720 278.430 297.685 ;
        RECT 279.550 295.720 284.410 297.685 ;
        RECT 285.530 295.720 290.390 297.685 ;
        RECT 291.510 295.720 296.370 297.685 ;
        RECT 2.860 4.280 297.060 295.720 ;
        RECT 2.860 2.050 20.830 4.280 ;
        RECT 21.950 2.050 63.610 4.280 ;
        RECT 64.730 2.050 106.390 4.280 ;
        RECT 107.510 2.050 149.170 4.280 ;
        RECT 150.290 2.050 191.950 4.280 ;
        RECT 193.070 2.050 234.730 4.280 ;
        RECT 235.850 2.050 277.510 4.280 ;
        RECT 278.630 2.050 297.060 4.280 ;
      LAYER met3 ;
        RECT 4.400 296.500 295.600 297.665 ;
        RECT 4.000 294.420 296.175 296.500 ;
        RECT 4.400 292.420 295.600 294.420 ;
        RECT 4.000 291.020 296.175 292.420 ;
        RECT 4.000 290.340 295.600 291.020 ;
        RECT 4.400 289.020 295.600 290.340 ;
        RECT 4.400 288.340 296.175 289.020 ;
        RECT 4.000 286.940 296.175 288.340 ;
        RECT 4.000 286.260 295.600 286.940 ;
        RECT 4.400 284.940 295.600 286.260 ;
        RECT 4.400 284.260 296.175 284.940 ;
        RECT 4.000 283.540 296.175 284.260 ;
        RECT 4.000 282.180 295.600 283.540 ;
        RECT 4.400 281.540 295.600 282.180 ;
        RECT 4.400 280.180 296.175 281.540 ;
        RECT 4.000 279.460 296.175 280.180 ;
        RECT 4.000 278.100 295.600 279.460 ;
        RECT 4.400 277.460 295.600 278.100 ;
        RECT 4.400 276.100 296.175 277.460 ;
        RECT 4.000 275.380 296.175 276.100 ;
        RECT 4.000 274.020 295.600 275.380 ;
        RECT 4.400 273.380 295.600 274.020 ;
        RECT 4.400 272.020 296.175 273.380 ;
        RECT 4.000 271.980 296.175 272.020 ;
        RECT 4.000 269.980 295.600 271.980 ;
        RECT 4.000 269.940 296.175 269.980 ;
        RECT 4.400 267.940 296.175 269.940 ;
        RECT 4.000 267.900 296.175 267.940 ;
        RECT 4.000 266.540 295.600 267.900 ;
        RECT 4.400 265.900 295.600 266.540 ;
        RECT 4.400 264.540 296.175 265.900 ;
        RECT 4.000 264.500 296.175 264.540 ;
        RECT 4.000 262.500 295.600 264.500 ;
        RECT 4.000 262.460 296.175 262.500 ;
        RECT 4.400 260.460 296.175 262.460 ;
        RECT 4.000 260.420 296.175 260.460 ;
        RECT 4.000 258.420 295.600 260.420 ;
        RECT 4.000 258.380 296.175 258.420 ;
        RECT 4.400 257.020 296.175 258.380 ;
        RECT 4.400 256.380 295.600 257.020 ;
        RECT 4.000 255.020 295.600 256.380 ;
        RECT 4.000 254.300 296.175 255.020 ;
        RECT 4.400 252.940 296.175 254.300 ;
        RECT 4.400 252.300 295.600 252.940 ;
        RECT 4.000 250.940 295.600 252.300 ;
        RECT 4.000 250.220 296.175 250.940 ;
        RECT 4.400 248.860 296.175 250.220 ;
        RECT 4.400 248.220 295.600 248.860 ;
        RECT 4.000 246.860 295.600 248.220 ;
        RECT 4.000 246.140 296.175 246.860 ;
        RECT 4.400 245.460 296.175 246.140 ;
        RECT 4.400 244.140 295.600 245.460 ;
        RECT 4.000 243.460 295.600 244.140 ;
        RECT 4.000 242.060 296.175 243.460 ;
        RECT 4.400 241.380 296.175 242.060 ;
        RECT 4.400 240.060 295.600 241.380 ;
        RECT 4.000 239.380 295.600 240.060 ;
        RECT 4.000 237.980 296.175 239.380 ;
        RECT 4.400 235.980 295.600 237.980 ;
        RECT 4.000 234.580 296.175 235.980 ;
        RECT 4.400 233.900 296.175 234.580 ;
        RECT 4.400 232.580 295.600 233.900 ;
        RECT 4.000 231.900 295.600 232.580 ;
        RECT 4.000 230.500 296.175 231.900 ;
        RECT 4.400 229.820 296.175 230.500 ;
        RECT 4.400 228.500 295.600 229.820 ;
        RECT 4.000 227.820 295.600 228.500 ;
        RECT 4.000 226.420 296.175 227.820 ;
        RECT 4.400 224.420 295.600 226.420 ;
        RECT 4.000 222.340 296.175 224.420 ;
        RECT 4.400 220.340 295.600 222.340 ;
        RECT 4.000 218.940 296.175 220.340 ;
        RECT 4.000 218.260 295.600 218.940 ;
        RECT 4.400 216.940 295.600 218.260 ;
        RECT 4.400 216.260 296.175 216.940 ;
        RECT 4.000 214.860 296.175 216.260 ;
        RECT 4.000 214.180 295.600 214.860 ;
        RECT 4.400 212.860 295.600 214.180 ;
        RECT 4.400 212.180 296.175 212.860 ;
        RECT 4.000 211.460 296.175 212.180 ;
        RECT 4.000 210.100 295.600 211.460 ;
        RECT 4.400 209.460 295.600 210.100 ;
        RECT 4.400 208.100 296.175 209.460 ;
        RECT 4.000 207.380 296.175 208.100 ;
        RECT 4.000 206.020 295.600 207.380 ;
        RECT 4.400 205.380 295.600 206.020 ;
        RECT 4.400 204.020 296.175 205.380 ;
        RECT 4.000 203.300 296.175 204.020 ;
        RECT 4.000 202.620 295.600 203.300 ;
        RECT 4.400 201.300 295.600 202.620 ;
        RECT 4.400 200.620 296.175 201.300 ;
        RECT 4.000 199.900 296.175 200.620 ;
        RECT 4.000 198.540 295.600 199.900 ;
        RECT 4.400 197.900 295.600 198.540 ;
        RECT 4.400 196.540 296.175 197.900 ;
        RECT 4.000 195.820 296.175 196.540 ;
        RECT 4.000 194.460 295.600 195.820 ;
        RECT 4.400 193.820 295.600 194.460 ;
        RECT 4.400 192.460 296.175 193.820 ;
        RECT 4.000 192.420 296.175 192.460 ;
        RECT 4.000 190.420 295.600 192.420 ;
        RECT 4.000 190.380 296.175 190.420 ;
        RECT 4.400 188.380 296.175 190.380 ;
        RECT 4.000 188.340 296.175 188.380 ;
        RECT 4.000 186.340 295.600 188.340 ;
        RECT 4.000 186.300 296.175 186.340 ;
        RECT 4.400 184.300 296.175 186.300 ;
        RECT 4.000 184.260 296.175 184.300 ;
        RECT 4.000 182.260 295.600 184.260 ;
        RECT 4.000 182.220 296.175 182.260 ;
        RECT 4.400 180.860 296.175 182.220 ;
        RECT 4.400 180.220 295.600 180.860 ;
        RECT 4.000 178.860 295.600 180.220 ;
        RECT 4.000 178.140 296.175 178.860 ;
        RECT 4.400 176.780 296.175 178.140 ;
        RECT 4.400 176.140 295.600 176.780 ;
        RECT 4.000 174.780 295.600 176.140 ;
        RECT 4.000 174.060 296.175 174.780 ;
        RECT 4.400 173.380 296.175 174.060 ;
        RECT 4.400 172.060 295.600 173.380 ;
        RECT 4.000 171.380 295.600 172.060 ;
        RECT 4.000 169.980 296.175 171.380 ;
        RECT 4.400 169.300 296.175 169.980 ;
        RECT 4.400 167.980 295.600 169.300 ;
        RECT 4.000 167.300 295.600 167.980 ;
        RECT 4.000 166.580 296.175 167.300 ;
        RECT 4.400 165.900 296.175 166.580 ;
        RECT 4.400 164.580 295.600 165.900 ;
        RECT 4.000 163.900 295.600 164.580 ;
        RECT 4.000 162.500 296.175 163.900 ;
        RECT 4.400 161.820 296.175 162.500 ;
        RECT 4.400 160.500 295.600 161.820 ;
        RECT 4.000 159.820 295.600 160.500 ;
        RECT 4.000 158.420 296.175 159.820 ;
        RECT 4.400 157.740 296.175 158.420 ;
        RECT 4.400 156.420 295.600 157.740 ;
        RECT 4.000 155.740 295.600 156.420 ;
        RECT 4.000 154.340 296.175 155.740 ;
        RECT 4.400 152.340 295.600 154.340 ;
        RECT 4.000 150.260 296.175 152.340 ;
        RECT 4.400 148.260 295.600 150.260 ;
        RECT 4.000 146.860 296.175 148.260 ;
        RECT 4.000 146.180 295.600 146.860 ;
        RECT 4.400 144.860 295.600 146.180 ;
        RECT 4.400 144.180 296.175 144.860 ;
        RECT 4.000 142.780 296.175 144.180 ;
        RECT 4.000 142.100 295.600 142.780 ;
        RECT 4.400 140.780 295.600 142.100 ;
        RECT 4.400 140.100 296.175 140.780 ;
        RECT 4.000 138.700 296.175 140.100 ;
        RECT 4.000 138.020 295.600 138.700 ;
        RECT 4.400 136.700 295.600 138.020 ;
        RECT 4.400 136.020 296.175 136.700 ;
        RECT 4.000 135.300 296.175 136.020 ;
        RECT 4.000 134.620 295.600 135.300 ;
        RECT 4.400 133.300 295.600 134.620 ;
        RECT 4.400 132.620 296.175 133.300 ;
        RECT 4.000 131.220 296.175 132.620 ;
        RECT 4.000 130.540 295.600 131.220 ;
        RECT 4.400 129.220 295.600 130.540 ;
        RECT 4.400 128.540 296.175 129.220 ;
        RECT 4.000 127.820 296.175 128.540 ;
        RECT 4.000 126.460 295.600 127.820 ;
        RECT 4.400 125.820 295.600 126.460 ;
        RECT 4.400 124.460 296.175 125.820 ;
        RECT 4.000 123.740 296.175 124.460 ;
        RECT 4.000 122.380 295.600 123.740 ;
        RECT 4.400 121.740 295.600 122.380 ;
        RECT 4.400 120.380 296.175 121.740 ;
        RECT 4.000 120.340 296.175 120.380 ;
        RECT 4.000 118.340 295.600 120.340 ;
        RECT 4.000 118.300 296.175 118.340 ;
        RECT 4.400 116.300 296.175 118.300 ;
        RECT 4.000 116.260 296.175 116.300 ;
        RECT 4.000 114.260 295.600 116.260 ;
        RECT 4.000 114.220 296.175 114.260 ;
        RECT 4.400 112.220 296.175 114.220 ;
        RECT 4.000 112.180 296.175 112.220 ;
        RECT 4.000 110.180 295.600 112.180 ;
        RECT 4.000 110.140 296.175 110.180 ;
        RECT 4.400 108.780 296.175 110.140 ;
        RECT 4.400 108.140 295.600 108.780 ;
        RECT 4.000 106.780 295.600 108.140 ;
        RECT 4.000 106.060 296.175 106.780 ;
        RECT 4.400 104.700 296.175 106.060 ;
        RECT 4.400 104.060 295.600 104.700 ;
        RECT 4.000 102.700 295.600 104.060 ;
        RECT 4.000 102.660 296.175 102.700 ;
        RECT 4.400 101.300 296.175 102.660 ;
        RECT 4.400 100.660 295.600 101.300 ;
        RECT 4.000 99.300 295.600 100.660 ;
        RECT 4.000 98.580 296.175 99.300 ;
        RECT 4.400 97.220 296.175 98.580 ;
        RECT 4.400 96.580 295.600 97.220 ;
        RECT 4.000 95.220 295.600 96.580 ;
        RECT 4.000 94.500 296.175 95.220 ;
        RECT 4.400 93.140 296.175 94.500 ;
        RECT 4.400 92.500 295.600 93.140 ;
        RECT 4.000 91.140 295.600 92.500 ;
        RECT 4.000 90.420 296.175 91.140 ;
        RECT 4.400 89.740 296.175 90.420 ;
        RECT 4.400 88.420 295.600 89.740 ;
        RECT 4.000 87.740 295.600 88.420 ;
        RECT 4.000 86.340 296.175 87.740 ;
        RECT 4.400 85.660 296.175 86.340 ;
        RECT 4.400 84.340 295.600 85.660 ;
        RECT 4.000 83.660 295.600 84.340 ;
        RECT 4.000 82.260 296.175 83.660 ;
        RECT 4.400 80.260 295.600 82.260 ;
        RECT 4.000 78.180 296.175 80.260 ;
        RECT 4.400 76.180 295.600 78.180 ;
        RECT 4.000 74.780 296.175 76.180 ;
        RECT 4.000 74.100 295.600 74.780 ;
        RECT 4.400 72.780 295.600 74.100 ;
        RECT 4.400 72.100 296.175 72.780 ;
        RECT 4.000 70.700 296.175 72.100 ;
        RECT 4.000 70.020 295.600 70.700 ;
        RECT 4.400 68.700 295.600 70.020 ;
        RECT 4.400 68.020 296.175 68.700 ;
        RECT 4.000 66.620 296.175 68.020 ;
        RECT 4.400 64.620 295.600 66.620 ;
        RECT 4.000 63.220 296.175 64.620 ;
        RECT 4.000 62.540 295.600 63.220 ;
        RECT 4.400 61.220 295.600 62.540 ;
        RECT 4.400 60.540 296.175 61.220 ;
        RECT 4.000 59.140 296.175 60.540 ;
        RECT 4.000 58.460 295.600 59.140 ;
        RECT 4.400 57.140 295.600 58.460 ;
        RECT 4.400 56.460 296.175 57.140 ;
        RECT 4.000 55.740 296.175 56.460 ;
        RECT 4.000 54.380 295.600 55.740 ;
        RECT 4.400 53.740 295.600 54.380 ;
        RECT 4.400 52.380 296.175 53.740 ;
        RECT 4.000 51.660 296.175 52.380 ;
        RECT 4.000 50.300 295.600 51.660 ;
        RECT 4.400 49.660 295.600 50.300 ;
        RECT 4.400 48.300 296.175 49.660 ;
        RECT 4.000 47.580 296.175 48.300 ;
        RECT 4.000 46.220 295.600 47.580 ;
        RECT 4.400 45.580 295.600 46.220 ;
        RECT 4.400 44.220 296.175 45.580 ;
        RECT 4.000 44.180 296.175 44.220 ;
        RECT 4.000 42.180 295.600 44.180 ;
        RECT 4.000 42.140 296.175 42.180 ;
        RECT 4.400 40.140 296.175 42.140 ;
        RECT 4.000 40.100 296.175 40.140 ;
        RECT 4.000 38.100 295.600 40.100 ;
        RECT 4.000 38.060 296.175 38.100 ;
        RECT 4.400 36.700 296.175 38.060 ;
        RECT 4.400 36.060 295.600 36.700 ;
        RECT 4.000 34.700 295.600 36.060 ;
        RECT 4.000 34.660 296.175 34.700 ;
        RECT 4.400 32.660 296.175 34.660 ;
        RECT 4.000 32.620 296.175 32.660 ;
        RECT 4.000 30.620 295.600 32.620 ;
        RECT 4.000 30.580 296.175 30.620 ;
        RECT 4.400 29.220 296.175 30.580 ;
        RECT 4.400 28.580 295.600 29.220 ;
        RECT 4.000 27.220 295.600 28.580 ;
        RECT 4.000 26.500 296.175 27.220 ;
        RECT 4.400 25.140 296.175 26.500 ;
        RECT 4.400 24.500 295.600 25.140 ;
        RECT 4.000 23.140 295.600 24.500 ;
        RECT 4.000 22.420 296.175 23.140 ;
        RECT 4.400 21.060 296.175 22.420 ;
        RECT 4.400 20.420 295.600 21.060 ;
        RECT 4.000 19.060 295.600 20.420 ;
        RECT 4.000 18.340 296.175 19.060 ;
        RECT 4.400 17.660 296.175 18.340 ;
        RECT 4.400 16.340 295.600 17.660 ;
        RECT 4.000 15.660 295.600 16.340 ;
        RECT 4.000 14.260 296.175 15.660 ;
        RECT 4.400 13.580 296.175 14.260 ;
        RECT 4.400 12.260 295.600 13.580 ;
        RECT 4.000 11.580 295.600 12.260 ;
        RECT 4.000 10.180 296.175 11.580 ;
        RECT 4.400 8.180 295.600 10.180 ;
        RECT 4.000 6.100 296.175 8.180 ;
        RECT 4.400 4.100 295.600 6.100 ;
        RECT 4.000 2.700 296.175 4.100 ;
        RECT 4.400 2.555 295.600 2.700 ;
      LAYER met4 ;
        RECT 95.975 17.175 97.440 271.825 ;
        RECT 99.840 17.175 174.240 271.825 ;
        RECT 176.640 17.175 251.040 271.825 ;
        RECT 253.440 17.175 288.585 271.825 ;
  END
END wrapped_vgademo_on_fpga
END LIBRARY

