* NGSPICE file created from wrapped_vgademo_on_fpga.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_8 abstract view
.subckt sky130_fd_sc_hd__ebufn_8 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_2 abstract view
.subckt sky130_fd_sc_hd__o32ai_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_4 abstract view
.subckt sky130_fd_sc_hd__or2b_4 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_4 abstract view
.subckt sky130_fd_sc_hd__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_2 abstract view
.subckt sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_1 abstract view
.subckt sky130_fd_sc_hd__o311ai_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

.subckt wrapped_vgademo_on_fpga active io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21]
+ io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29]
+ io_in[2] io_in[30] io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37]
+ io_in[3] io_in[4] io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10]
+ io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18]
+ io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25]
+ io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32]
+ io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5]
+ io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12]
+ io_out[13] io_out[14] io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1]
+ io_out[20] io_out[21] io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27]
+ io_out[28] io_out[29] io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34]
+ io_out[35] io_out[36] io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ io_out[8] io_out[9] la1_data_in[0] la1_data_in[10] la1_data_in[11] la1_data_in[12]
+ la1_data_in[13] la1_data_in[14] la1_data_in[15] la1_data_in[16] la1_data_in[17]
+ la1_data_in[18] la1_data_in[19] la1_data_in[1] la1_data_in[20] la1_data_in[21] la1_data_in[22]
+ la1_data_in[23] la1_data_in[24] la1_data_in[25] la1_data_in[26] la1_data_in[27]
+ la1_data_in[28] la1_data_in[29] la1_data_in[2] la1_data_in[30] la1_data_in[31] la1_data_in[3]
+ la1_data_in[4] la1_data_in[5] la1_data_in[6] la1_data_in[7] la1_data_in[8] la1_data_in[9]
+ la1_data_out[0] la1_data_out[10] la1_data_out[11] la1_data_out[12] la1_data_out[13]
+ la1_data_out[14] la1_data_out[15] la1_data_out[16] la1_data_out[17] la1_data_out[18]
+ la1_data_out[19] la1_data_out[1] la1_data_out[20] la1_data_out[21] la1_data_out[22]
+ la1_data_out[23] la1_data_out[24] la1_data_out[25] la1_data_out[26] la1_data_out[27]
+ la1_data_out[28] la1_data_out[29] la1_data_out[2] la1_data_out[30] la1_data_out[31]
+ la1_data_out[3] la1_data_out[4] la1_data_out[5] la1_data_out[6] la1_data_out[7]
+ la1_data_out[8] la1_data_out[9] la1_oenb[0] la1_oenb[10] la1_oenb[11] la1_oenb[12]
+ la1_oenb[13] la1_oenb[14] la1_oenb[15] la1_oenb[16] la1_oenb[17] la1_oenb[18] la1_oenb[19]
+ la1_oenb[1] la1_oenb[20] la1_oenb[21] la1_oenb[22] la1_oenb[23] la1_oenb[24] la1_oenb[25]
+ la1_oenb[26] la1_oenb[27] la1_oenb[28] la1_oenb[29] la1_oenb[2] la1_oenb[30] la1_oenb[31]
+ la1_oenb[3] la1_oenb[4] la1_oenb[5] la1_oenb[6] la1_oenb[7] la1_oenb[8] la1_oenb[9]
+ vccd1 vssd1 wb_clk_i
XFILLER_79_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7963_ _7963_/A vssd1 vssd1 vccd1 vccd1 _8134_/B sky130_fd_sc_hd__buf_2
XFILLER_82_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6914_ _6914_/A _6914_/B _6914_/C vssd1 vssd1 vccd1 vccd1 _7044_/A sky130_fd_sc_hd__and3_1
XFILLER_54_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7894_ _7894_/A _7894_/B _7894_/C vssd1 vssd1 vccd1 vccd1 _7949_/B sky130_fd_sc_hd__nand3_1
X_6845_ _7107_/A _7443_/A vssd1 vssd1 vccd1 vccd1 _7088_/A sky130_fd_sc_hd__nand2_1
XFILLER_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6776_ _8703_/Q vssd1 vssd1 vccd1 vccd1 _7533_/A sky130_fd_sc_hd__inv_2
X_8515_ _7503_/X _8715_/Q _8510_/X _8514_/X vssd1 vssd1 vccd1 vccd1 _8715_/D sky130_fd_sc_hd__o22a_1
X_5727_ _5731_/A _5727_/B vssd1 vssd1 vccd1 vccd1 _5792_/B sky130_fd_sc_hd__xor2_2
X_8446_ _8382_/A _8308_/A _8446_/S vssd1 vssd1 vccd1 vccd1 _8447_/B sky130_fd_sc_hd__mux2_1
X_5658_ _5658_/A vssd1 vssd1 vccd1 vccd1 _5922_/A sky130_fd_sc_hd__clkbuf_2
X_8377_ _8377_/A _8377_/B vssd1 vssd1 vccd1 vccd1 _8377_/Y sky130_fd_sc_hd__nor2_1
X_4609_ _8578_/Q _4610_/C _4608_/Y vssd1 vssd1 vccd1 vccd1 _8578_/D sky130_fd_sc_hd__a21oi_1
X_5589_ _5589_/A _5589_/B vssd1 vssd1 vccd1 vccd1 _5590_/B sky130_fd_sc_hd__xor2_1
X_7328_ _7373_/A _7373_/B vssd1 vssd1 vccd1 vccd1 _7330_/B sky130_fd_sc_hd__and2_1
XFILLER_104_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7259_ _7259_/A _7259_/B vssd1 vssd1 vccd1 vccd1 _7260_/B sky130_fd_sc_hd__and2_1
XFILLER_89_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4960_ _4960_/A _4961_/B vssd1 vssd1 vccd1 vccd1 _5054_/C sky130_fd_sc_hd__nor2_2
XFILLER_17_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4891_ _4922_/A vssd1 vssd1 vccd1 vccd1 _5243_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6630_ _6614_/X _6657_/B _6657_/C _6798_/A _7245_/A vssd1 vssd1 vccd1 vccd1 _6639_/A
+ sky130_fd_sc_hd__a311o_1
X_6561_ _6561_/A _6561_/B vssd1 vssd1 vccd1 vccd1 _6562_/B sky130_fd_sc_hd__nor2_2
X_8300_ _8241_/A _8241_/B _8299_/X vssd1 vssd1 vccd1 vccd1 _8346_/A sky130_fd_sc_hd__a21oi_1
X_5512_ _5512_/A _5560_/B vssd1 vssd1 vccd1 vccd1 _5513_/B sky130_fd_sc_hd__xnor2_1
X_6492_ _6481_/Y _6491_/X _4784_/A vssd1 vssd1 vccd1 vccd1 _8686_/D sky130_fd_sc_hd__a21oi_1
X_8231_ _8232_/A _8410_/B vssd1 vssd1 vccd1 vccd1 _8337_/B sky130_fd_sc_hd__or2_1
XFILLER_8_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5443_ _5442_/A _5442_/B _5442_/C _5447_/B vssd1 vssd1 vccd1 vccd1 _5444_/B sky130_fd_sc_hd__a22oi_1
X_8162_ _8254_/B _8162_/B vssd1 vssd1 vccd1 vccd1 _8163_/B sky130_fd_sc_hd__nor2_1
X_5374_ _5374_/A _5374_/B _5374_/C vssd1 vssd1 vccd1 vccd1 _5375_/A sky130_fd_sc_hd__and3_1
X_7113_ _7113_/A _7113_/B vssd1 vssd1 vccd1 vccd1 _7123_/A sky130_fd_sc_hd__xnor2_1
X_8093_ _8097_/A _8097_/B _8093_/C _8093_/D vssd1 vssd1 vccd1 vccd1 _8500_/B sky130_fd_sc_hd__and4bb_1
XFILLER_86_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7044_ _7044_/A _7044_/B _7044_/C _7044_/D vssd1 vssd1 vccd1 vccd1 _7044_/X sky130_fd_sc_hd__or4_2
XFILLER_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7946_ _8097_/B _7946_/B vssd1 vssd1 vccd1 vccd1 _7946_/X sky130_fd_sc_hd__xor2_2
XFILLER_55_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7877_ _7877_/A _8406_/A vssd1 vssd1 vccd1 vccd1 _7877_/Y sky130_fd_sc_hd__nor2_1
XFILLER_42_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6828_ _6647_/A _7265_/A _6730_/B _6827_/X vssd1 vssd1 vccd1 vccd1 _6850_/A sky130_fd_sc_hd__o31a_2
XFILLER_11_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6759_ _7185_/A _6756_/X _6757_/Y _6758_/X vssd1 vssd1 vccd1 vccd1 _6787_/A sky130_fd_sc_hd__a31o_1
XFILLER_10_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8429_ _8429_/A _8429_/B vssd1 vssd1 vccd1 vccd1 _8431_/B sky130_fd_sc_hd__xnor2_1
XFILLER_12_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8745__23 vssd1 vssd1 vccd1 vccd1 _8745__23/HI _8840_/A sky130_fd_sc_hd__conb_1
XFILLER_61_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5090_ _5231_/A _5084_/X _5252_/B _5088_/X _5089_/Y vssd1 vssd1 vccd1 vccd1 _5090_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_83_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7800_ _7800_/A _7800_/B vssd1 vssd1 vccd1 vccd1 _7801_/B sky130_fd_sc_hd__xnor2_1
XFILLER_52_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5992_ _5990_/A _5888_/B _5916_/B _5915_/B _5915_/A vssd1 vssd1 vccd1 vccd1 _6199_/A
+ sky130_fd_sc_hd__a32o_1
XFILLER_91_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7731_ _7746_/A vssd1 vssd1 vccd1 vccd1 _8205_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_52_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4943_ _5098_/D _5153_/B vssd1 vssd1 vccd1 vccd1 _5172_/C sky130_fd_sc_hd__or2_1
X_7662_ _7664_/A _7995_/B vssd1 vssd1 vccd1 vccd1 _7666_/C sky130_fd_sc_hd__nor2_1
XFILLER_60_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6613_ _6628_/A _8611_/Q vssd1 vssd1 vccd1 vccd1 _6656_/B sky130_fd_sc_hd__or2_1
X_4874_ _5010_/B _4898_/B vssd1 vssd1 vccd1 vccd1 _5006_/A sky130_fd_sc_hd__nor2_1
X_7593_ _8707_/Q _7593_/B vssd1 vssd1 vccd1 vccd1 _7594_/B sky130_fd_sc_hd__and2b_1
XFILLER_20_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6544_ _8694_/Q vssd1 vssd1 vccd1 vccd1 _6628_/A sky130_fd_sc_hd__inv_2
X_6475_ _8629_/Q _6475_/B _8633_/Q _6475_/D vssd1 vssd1 vccd1 vccd1 _6477_/B sky130_fd_sc_hd__or4_1
X_8214_ _8214_/A _8214_/B vssd1 vssd1 vccd1 vccd1 _8214_/Y sky130_fd_sc_hd__nand2_1
X_5426_ _5424_/Y _5425_/X _5419_/X vssd1 vssd1 vccd1 vccd1 _5426_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_87_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8145_ _8196_/A _8361_/A _8144_/Y vssd1 vssd1 vccd1 vccd1 _8146_/B sky130_fd_sc_hd__o21bai_2
X_5357_ _6511_/A vssd1 vssd1 vccd1 vccd1 _5357_/X sky130_fd_sc_hd__clkbuf_2
XINSDIODE2_4 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8076_ _8305_/A vssd1 vssd1 vccd1 vccd1 _8141_/A sky130_fd_sc_hd__inv_2
X_5288_ _8618_/Q _5288_/B vssd1 vssd1 vccd1 vccd1 _5288_/X sky130_fd_sc_hd__or2_1
XFILLER_101_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7027_ _7027_/A _7027_/B vssd1 vssd1 vccd1 vccd1 _7036_/A sky130_fd_sc_hd__xnor2_1
XFILLER_75_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7929_ _7929_/A _7929_/B _7929_/C vssd1 vssd1 vccd1 vccd1 _7929_/X sky130_fd_sc_hd__and3_1
XFILLER_70_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4590_ _8572_/Q _8571_/Q _8573_/Q vssd1 vssd1 vccd1 vccd1 _4591_/C sky130_fd_sc_hd__a21o_1
X_6260_ _6260_/A _6260_/B vssd1 vssd1 vccd1 vccd1 _6261_/B sky130_fd_sc_hd__xnor2_1
X_6191_ _5969_/A _5969_/B _6190_/X vssd1 vssd1 vccd1 vccd1 _6192_/B sky130_fd_sc_hd__a21oi_1
X_5211_ _5226_/B _5127_/A _4786_/B vssd1 vssd1 vccd1 vccd1 _5212_/S sky130_fd_sc_hd__o21a_1
X_5142_ _5253_/A _5139_/X _5132_/X _4661_/A _5141_/X vssd1 vssd1 vccd1 vccd1 _5142_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_96_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5073_ _5231_/A _5145_/B _5071_/X _5072_/X _4686_/A vssd1 vssd1 vccd1 vccd1 _5073_/X
+ sky130_fd_sc_hd__o41a_1
X_8901_ _8901_/A _4418_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[10] sky130_fd_sc_hd__ebufn_8
XFILLER_92_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8832_ _8832_/A _4342_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[11] sky130_fd_sc_hd__ebufn_8
XFILLER_80_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5975_ _5975_/A _6173_/B vssd1 vssd1 vccd1 vccd1 _5976_/B sky130_fd_sc_hd__xnor2_1
X_7714_ _7722_/A _7714_/B vssd1 vssd1 vccd1 vccd1 _7887_/A sky130_fd_sc_hd__and2_2
X_4926_ _5193_/B _5057_/C vssd1 vssd1 vccd1 vccd1 _4939_/A sky130_fd_sc_hd__or2_1
X_8694_ input3/X _8694_/D vssd1 vssd1 vccd1 vccd1 _8694_/Q sky130_fd_sc_hd__dfxtp_1
X_7645_ _7986_/A _7796_/A vssd1 vssd1 vccd1 vccd1 _7682_/A sky130_fd_sc_hd__nand2_2
X_4857_ _5041_/A _4857_/B vssd1 vssd1 vccd1 vccd1 _5116_/B sky130_fd_sc_hd__nor2_1
XFILLER_33_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7576_ _7593_/B _7587_/A _7604_/A vssd1 vssd1 vccd1 vccd1 _7576_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4788_ _4864_/B vssd1 vssd1 vccd1 vccd1 _4903_/A sky130_fd_sc_hd__inv_2
X_6527_ _6525_/Y _6527_/B vssd1 vssd1 vccd1 vccd1 _6529_/A sky130_fd_sc_hd__and2b_1
XFILLER_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6458_ _6459_/B _6459_/C _6457_/Y vssd1 vssd1 vccd1 vccd1 _8681_/D sky130_fd_sc_hd__a21oi_1
XFILLER_69_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5409_ _8647_/Q vssd1 vssd1 vccd1 vccd1 _5607_/A sky130_fd_sc_hd__inv_2
X_6389_ _8678_/Q vssd1 vssd1 vccd1 vccd1 _6450_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_102_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8128_ _8128_/A _8205_/C vssd1 vssd1 vccd1 vccd1 _8130_/B sky130_fd_sc_hd__xnor2_1
XFILLER_87_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8059_ _8172_/A _8058_/X vssd1 vssd1 vccd1 vccd1 _8140_/A sky130_fd_sc_hd__or2b_1
XFILLER_55_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5760_ _6123_/A _5674_/A _5974_/A vssd1 vssd1 vccd1 vccd1 _5777_/B sky130_fd_sc_hd__a21o_1
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5691_ _6044_/A _6180_/A vssd1 vssd1 vccd1 vccd1 _5692_/B sky130_fd_sc_hd__nor2_1
XFILLER_30_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4711_ _4739_/A _4681_/B _5127_/A _5226_/B vssd1 vssd1 vccd1 vccd1 _4712_/C sky130_fd_sc_hd__a31o_1
X_7430_ _7449_/A _7449_/B _7449_/C vssd1 vssd1 vccd1 vccd1 _7473_/B sky130_fd_sc_hd__a21o_1
X_4642_ _8589_/Q _4641_/B _4607_/X vssd1 vssd1 vccd1 vccd1 _4643_/B sky130_fd_sc_hd__o21ai_1
X_7361_ _7354_/A _7354_/B _7360_/X vssd1 vssd1 vccd1 vccd1 _7454_/A sky130_fd_sc_hd__o21ba_1
X_4573_ _8578_/Q _8577_/Q _8580_/Q _4573_/D vssd1 vssd1 vccd1 vccd1 _4579_/B sky130_fd_sc_hd__or4_1
X_7292_ _7377_/A _7377_/B vssd1 vssd1 vccd1 vccd1 _7332_/A sky130_fd_sc_hd__nor2_1
X_6312_ _6312_/A _6312_/B vssd1 vssd1 vccd1 vccd1 _6314_/A sky130_fd_sc_hd__nand2_1
XFILLER_103_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6243_ _6244_/A _6243_/B vssd1 vssd1 vccd1 vccd1 _6317_/B sky130_fd_sc_hd__xnor2_2
X_6174_ _5976_/A _5976_/B _6173_/X vssd1 vssd1 vccd1 vccd1 _6241_/A sky130_fd_sc_hd__a21oi_2
XFILLER_69_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5125_ _5125_/A _5248_/A _4952_/A vssd1 vssd1 vccd1 vccd1 _5125_/X sky130_fd_sc_hd__or3b_1
X_5056_ _5214_/C _5098_/D _5053_/X _5055_/X vssd1 vssd1 vccd1 vccd1 _5057_/D sky130_fd_sc_hd__o31a_1
XFILLER_29_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5958_ _5958_/A vssd1 vssd1 vccd1 vccd1 _6183_/A sky130_fd_sc_hd__clkbuf_2
X_4909_ _4909_/A _5011_/A _5026_/B vssd1 vssd1 vccd1 vccd1 _4975_/B sky130_fd_sc_hd__or3b_1
X_8677_ input3/X _8677_/D vssd1 vssd1 vccd1 vccd1 _8677_/Q sky130_fd_sc_hd__dfxtp_1
X_5889_ _5890_/B _5889_/B vssd1 vssd1 vccd1 vccd1 _5889_/X sky130_fd_sc_hd__and2b_1
X_7628_ _7673_/A _7673_/B vssd1 vssd1 vccd1 vccd1 _7664_/A sky130_fd_sc_hd__nor2_2
XFILLER_21_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7559_ _8539_/A _8531_/A _8719_/Q _8552_/B _8546_/A vssd1 vssd1 vccd1 vccd1 _7559_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_20_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6930_ _7065_/A _7065_/B vssd1 vssd1 vccd1 vccd1 _6931_/B sky130_fd_sc_hd__xor2_1
XFILLER_47_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6861_ _6869_/A _6864_/A vssd1 vssd1 vccd1 vccd1 _6862_/A sky130_fd_sc_hd__nor2_1
X_6792_ _6919_/B vssd1 vssd1 vccd1 vccd1 _7046_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_22_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8600_ input3/X _8600_/D vssd1 vssd1 vccd1 vccd1 _8600_/Q sky130_fd_sc_hd__dfxtp_2
X_5812_ _5812_/A _5812_/B vssd1 vssd1 vccd1 vccd1 _5813_/B sky130_fd_sc_hd__nor2_1
X_8531_ _8531_/A _8706_/Q vssd1 vssd1 vccd1 vccd1 _8533_/B sky130_fd_sc_hd__xor2_1
X_5743_ _5742_/A _5740_/Y _5920_/A vssd1 vssd1 vccd1 vccd1 _5744_/B sky130_fd_sc_hd__a21oi_1
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8462_ _8462_/A _8462_/B _8462_/C vssd1 vssd1 vccd1 vccd1 _8462_/Y sky130_fd_sc_hd__nor3_1
X_5674_ _5674_/A _6193_/A vssd1 vssd1 vccd1 vccd1 _5675_/B sky130_fd_sc_hd__xnor2_2
XFILLER_30_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8393_ _8333_/B _8393_/B vssd1 vssd1 vccd1 vccd1 _8400_/B sky130_fd_sc_hd__and2b_1
X_7413_ _7413_/A _7449_/A vssd1 vssd1 vccd1 vccd1 _7452_/B sky130_fd_sc_hd__and2_1
X_4625_ _4628_/C _4625_/B vssd1 vssd1 vccd1 vccd1 _8583_/D sky130_fd_sc_hd__nor2_1
X_4556_ _4556_/A vssd1 vssd1 vccd1 vccd1 _8875_/A sky130_fd_sc_hd__clkbuf_1
X_7344_ _7345_/A _7345_/B _7345_/C vssd1 vssd1 vccd1 vccd1 _7344_/Y sky130_fd_sc_hd__o21ai_1
X_7275_ _7275_/A _7275_/B vssd1 vssd1 vccd1 vccd1 _7353_/B sky130_fd_sc_hd__xnor2_1
X_4487_ _7658_/B vssd1 vssd1 vccd1 vccd1 _4775_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6226_ _6226_/A vssd1 vssd1 vccd1 vccd1 _6226_/Y sky130_fd_sc_hd__clkinv_2
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6157_ _6157_/A _6157_/B vssd1 vssd1 vccd1 vccd1 _6164_/D sky130_fd_sc_hd__xor2_2
XFILLER_97_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5108_ _5245_/A _5243_/B _5256_/A _4990_/Y _4969_/B vssd1 vssd1 vccd1 vccd1 _5111_/A
+ sky130_fd_sc_hd__o32a_1
X_6088_ _6094_/A _6088_/B vssd1 vssd1 vccd1 vccd1 _6134_/B sky130_fd_sc_hd__nand2_1
X_5039_ _4928_/A _5038_/Y _5245_/A vssd1 vssd1 vccd1 vccd1 _5040_/C sky130_fd_sc_hd__a21oi_1
XFILLER_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8790__68 vssd1 vssd1 vccd1 vccd1 _8790__68/HI _8899_/A sky130_fd_sc_hd__conb_1
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4410_ _4414_/A vssd1 vssd1 vccd1 vccd1 _4410_/Y sky130_fd_sc_hd__inv_2
X_5390_ _6371_/A _8662_/Q _5386_/X _5389_/Y _8536_/A vssd1 vssd1 vccd1 vccd1 _5391_/A
+ sky130_fd_sc_hd__o311a_1
XFILLER_99_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4341_ _4365_/A vssd1 vssd1 vccd1 vccd1 _4346_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_98_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7060_ _7060_/A _7060_/B _7060_/C vssd1 vssd1 vccd1 vccd1 _7101_/C sky130_fd_sc_hd__nand3_2
XFILLER_98_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6011_ _6012_/B _6011_/B vssd1 vssd1 vccd1 vccd1 _6013_/A sky130_fd_sc_hd__and2b_1
XFILLER_100_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7962_ _8218_/A _7962_/B vssd1 vssd1 vccd1 vccd1 _7966_/A sky130_fd_sc_hd__nand2_1
XFILLER_82_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6913_ _6728_/A _6801_/A _7135_/A _6803_/B vssd1 vssd1 vccd1 vccd1 _6914_/C sky130_fd_sc_hd__a22o_1
XFILLER_54_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7893_ _7980_/A _7893_/B vssd1 vssd1 vccd1 vccd1 _7894_/C sky130_fd_sc_hd__and2b_1
X_6844_ _6844_/A _7193_/A vssd1 vssd1 vccd1 vccd1 _7443_/A sky130_fd_sc_hd__nor2_4
XFILLER_50_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6775_ _6710_/A _6712_/A _6710_/B _6605_/X vssd1 vssd1 vccd1 vccd1 _6779_/A sky130_fd_sc_hd__a31o_1
XFILLER_50_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8514_ _7946_/X _8527_/B _8513_/Y _8557_/A vssd1 vssd1 vccd1 vccd1 _8514_/X sky130_fd_sc_hd__a31o_1
XFILLER_10_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5726_ _5726_/A _5809_/A vssd1 vssd1 vccd1 vccd1 _5727_/B sky130_fd_sc_hd__xor2_2
X_8445_ _8445_/A _8445_/B _8445_/C vssd1 vssd1 vccd1 vccd1 _8447_/A sky130_fd_sc_hd__and3_1
X_5657_ _5657_/A _5657_/B vssd1 vssd1 vccd1 vccd1 _5658_/A sky130_fd_sc_hd__xor2_1
X_8376_ _8376_/A vssd1 vssd1 vccd1 vccd1 _8376_/Y sky130_fd_sc_hd__inv_2
X_4608_ _8578_/Q _4610_/C _4607_/X vssd1 vssd1 vccd1 vccd1 _4608_/Y sky130_fd_sc_hd__o21ai_1
X_5588_ _6213_/A _5795_/A _5587_/Y vssd1 vssd1 vccd1 vccd1 _5589_/B sky130_fd_sc_hd__a21oi_1
XFILLER_89_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7327_ _7327_/A _7327_/B vssd1 vssd1 vccd1 vccd1 _7373_/B sky130_fd_sc_hd__xor2_1
X_4539_ _8604_/Q _8603_/Q _5607_/B vssd1 vssd1 vccd1 vccd1 _4822_/C sky130_fd_sc_hd__o21a_2
X_7258_ _7258_/A _7258_/B vssd1 vssd1 vccd1 vccd1 _7259_/B sky130_fd_sc_hd__or2_1
XFILLER_89_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6209_ _6209_/A _6209_/B vssd1 vssd1 vccd1 vccd1 _6237_/A sky130_fd_sc_hd__xnor2_1
X_7189_ _7272_/A _7272_/B _7188_/X vssd1 vssd1 vccd1 vccd1 _7191_/A sky130_fd_sc_hd__o21ai_1
XFILLER_58_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4890_ _4890_/A vssd1 vssd1 vccd1 vccd1 _5092_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_44_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6560_ _8701_/Q _6560_/B vssd1 vssd1 vccd1 vccd1 _6561_/B sky130_fd_sc_hd__and2b_1
X_5511_ _5511_/A _5563_/A vssd1 vssd1 vccd1 vccd1 _5560_/B sky130_fd_sc_hd__xnor2_1
XFILLER_8_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6491_ _6486_/X _6488_/X _7537_/A _7529_/A vssd1 vssd1 vccd1 vccd1 _6491_/X sky130_fd_sc_hd__a211o_1
X_8230_ _8230_/A _8230_/B vssd1 vssd1 vccd1 vccd1 _8410_/B sky130_fd_sc_hd__nor2_1
X_5442_ _5442_/A _5442_/B _5442_/C _5447_/B vssd1 vssd1 vccd1 vccd1 _5444_/A sky130_fd_sc_hd__and4_1
X_8161_ _8161_/A _8161_/B vssd1 vssd1 vccd1 vccd1 _8162_/B sky130_fd_sc_hd__nor2_1
X_5373_ _8642_/Q _5373_/B vssd1 vssd1 vccd1 vccd1 _5374_/C sky130_fd_sc_hd__nand2_1
XFILLER_99_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7112_ _7112_/A _7112_/B vssd1 vssd1 vccd1 vccd1 _7113_/B sky130_fd_sc_hd__xnor2_1
X_8092_ _8015_/B _8015_/C _8015_/A vssd1 vssd1 vccd1 vccd1 _8093_/D sky130_fd_sc_hd__a21o_1
X_7043_ _7044_/C vssd1 vssd1 vccd1 vccd1 _7043_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7945_ _8097_/A _8094_/A vssd1 vssd1 vccd1 vccd1 _7946_/B sky130_fd_sc_hd__nand2_1
X_7876_ _7752_/A _7751_/B _7752_/B _7875_/X _7823_/A vssd1 vssd1 vccd1 vccd1 _8406_/A
+ sky130_fd_sc_hd__o311a_2
XFILLER_35_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6827_ _6827_/A _6731_/B vssd1 vssd1 vccd1 vccd1 _6827_/X sky130_fd_sc_hd__or2b_1
XFILLER_23_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6758_ _7184_/A _7313_/A _7180_/A vssd1 vssd1 vccd1 vccd1 _6758_/X sky130_fd_sc_hd__and3b_1
XFILLER_10_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6689_ _6689_/A _6695_/A _7047_/A vssd1 vssd1 vccd1 vccd1 _6689_/X sky130_fd_sc_hd__and3_1
X_5709_ _5768_/B _5710_/B _5709_/C vssd1 vssd1 vccd1 vccd1 _5783_/A sky130_fd_sc_hd__and3_1
X_8428_ _8428_/A _8428_/B vssd1 vssd1 vccd1 vccd1 _8431_/A sky130_fd_sc_hd__or2_1
XFILLER_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8359_ _8310_/A _8310_/B _8384_/B _8382_/A vssd1 vssd1 vccd1 vccd1 _8441_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_2_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8760__38 vssd1 vssd1 vccd1 vccd1 _8760__38/HI _8855_/A sky130_fd_sc_hd__conb_1
XFILLER_68_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5991_ _5991_/A _5991_/B vssd1 vssd1 vccd1 vccd1 _6198_/A sky130_fd_sc_hd__xnor2_2
X_7730_ _7814_/A _7814_/B vssd1 vssd1 vccd1 vccd1 _7815_/A sky130_fd_sc_hd__or2_1
XFILLER_64_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4942_ _4920_/X _4928_/Y _4941_/X _4970_/A vssd1 vssd1 vccd1 vccd1 _4942_/X sky130_fd_sc_hd__o211a_1
X_7661_ _8305_/A vssd1 vssd1 vccd1 vccd1 _7995_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6612_ _6751_/A vssd1 vssd1 vccd1 vccd1 _7219_/A sky130_fd_sc_hd__clkbuf_2
X_4873_ _5026_/B _5026_/C vssd1 vssd1 vccd1 vccd1 _5104_/B sky130_fd_sc_hd__and2_1
XFILLER_32_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7592_ _7592_/A vssd1 vssd1 vccd1 vccd1 _8709_/D sky130_fd_sc_hd__clkbuf_1
X_6543_ _6513_/X _6542_/X _6539_/A _7533_/B vssd1 vssd1 vccd1 vccd1 _8693_/D sky130_fd_sc_hd__o2bb2a_1
X_6474_ _8627_/Q _8626_/Q vssd1 vssd1 vccd1 vccd1 _6477_/A sky130_fd_sc_hd__nand2_1
X_8213_ _8312_/A _8213_/B vssd1 vssd1 vccd1 vccd1 _8239_/A sky130_fd_sc_hd__and2_2
X_5425_ _5425_/A _5425_/B vssd1 vssd1 vccd1 vccd1 _5425_/X sky130_fd_sc_hd__and2_1
X_8144_ _8147_/A _8060_/B _8305_/B vssd1 vssd1 vccd1 vccd1 _8144_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5356_ _8637_/Q _5360_/C vssd1 vssd1 vccd1 vccd1 _5359_/A sky130_fd_sc_hd__and2_1
XFILLER_101_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8075_ _7836_/B _8446_/S _8296_/A vssd1 vssd1 vccd1 vccd1 _8079_/A sky130_fd_sc_hd__o21ai_1
XINSDIODE2_5 _8527_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5287_ _8716_/Q _5285_/X _5286_/X _5283_/X vssd1 vssd1 vccd1 vccd1 _8617_/D sky130_fd_sc_hd__o211a_1
X_7026_ _6950_/A _6950_/B _7025_/X vssd1 vssd1 vccd1 vccd1 _7027_/B sky130_fd_sc_hd__a21oi_1
XFILLER_74_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7928_ _8018_/A _7928_/B vssd1 vssd1 vccd1 vccd1 _7929_/C sky130_fd_sc_hd__nor2_1
XFILLER_55_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7859_ _8395_/A _8116_/C vssd1 vssd1 vccd1 vccd1 _7859_/Y sky130_fd_sc_hd__nor2_1
XFILLER_11_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8805__83 vssd1 vssd1 vccd1 vccd1 _8805__83/HI _8914_/A sky130_fd_sc_hd__conb_1
XFILLER_93_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5210_ _5261_/A _5148_/X _5161_/X _5209_/X vssd1 vssd1 vccd1 vccd1 _5210_/X sky130_fd_sc_hd__o31a_1
X_6190_ _5970_/B _6190_/B vssd1 vssd1 vccd1 vccd1 _6190_/X sky130_fd_sc_hd__and2b_1
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5141_ _5224_/C _5133_/Y _5159_/C _5137_/X _5094_/B vssd1 vssd1 vccd1 vccd1 _5141_/X
+ sky130_fd_sc_hd__o32a_1
X_5072_ _5174_/B _5072_/B _5072_/C vssd1 vssd1 vccd1 vccd1 _5072_/X sky130_fd_sc_hd__or3_1
XFILLER_96_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8900_ _8900_/A _4416_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[9] sky130_fd_sc_hd__ebufn_8
XFILLER_56_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8831_ _8831_/A _4339_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[10] sky130_fd_sc_hd__ebufn_8
XFILLER_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7713_ _7886_/A vssd1 vssd1 vccd1 vccd1 _7853_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_5974_ _5974_/A _5974_/B vssd1 vssd1 vccd1 vccd1 _6173_/B sky130_fd_sc_hd__xnor2_1
X_4925_ _5116_/B _5241_/B vssd1 vssd1 vccd1 vccd1 _5057_/C sky130_fd_sc_hd__or2_2
X_8693_ input3/X _8693_/D vssd1 vssd1 vccd1 vccd1 _8693_/Q sky130_fd_sc_hd__dfxtp_1
X_7644_ _7644_/A _7644_/B vssd1 vssd1 vccd1 vccd1 _7796_/A sky130_fd_sc_hd__nor2_1
X_4856_ _4856_/A _5041_/A vssd1 vssd1 vccd1 vccd1 _5202_/A sky130_fd_sc_hd__nor2_2
X_7575_ _7616_/A _7571_/Y _7611_/A _7574_/X vssd1 vssd1 vccd1 vccd1 _7575_/Y sky130_fd_sc_hd__a31oi_1
X_6526_ _6526_/A _6526_/B vssd1 vssd1 vccd1 vccd1 _6527_/B sky130_fd_sc_hd__nand2_1
X_4787_ _4831_/C _4787_/B vssd1 vssd1 vccd1 vccd1 _4864_/B sky130_fd_sc_hd__nor2_1
XFILLER_20_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6457_ _6459_/B _6459_/C _6419_/X vssd1 vssd1 vccd1 vccd1 _6457_/Y sky130_fd_sc_hd__o21ai_1
X_6388_ _6441_/B _8673_/Q _6386_/X _6387_/X vssd1 vssd1 vccd1 vccd1 _6388_/X sky130_fd_sc_hd__a31o_1
X_5408_ _6507_/A _5449_/B vssd1 vssd1 vccd1 vccd1 _5413_/A sky130_fd_sc_hd__nor2_2
X_8127_ _8127_/A _8127_/B vssd1 vssd1 vccd1 vccd1 _8205_/C sky130_fd_sc_hd__xor2_1
X_5339_ _5342_/C _5339_/B vssd1 vssd1 vccd1 vccd1 _8631_/D sky130_fd_sc_hd__nor2_1
XFILLER_102_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8058_ _8057_/A _8280_/A _8057_/D _8057_/C vssd1 vssd1 vccd1 vccd1 _8058_/X sky130_fd_sc_hd__a31o_1
XFILLER_47_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7009_ _7010_/A _7010_/B _7010_/C vssd1 vssd1 vccd1 vccd1 _7011_/A sky130_fd_sc_hd__a21o_1
XFILLER_90_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5690_ _5961_/A _5961_/B vssd1 vssd1 vccd1 vccd1 _6107_/B sky130_fd_sc_hd__nand2_2
X_4710_ _4710_/A _4786_/B vssd1 vssd1 vccd1 vccd1 _4716_/B sky130_fd_sc_hd__nor2_1
X_4641_ _8589_/Q _4641_/B vssd1 vssd1 vccd1 vccd1 _4645_/B sky130_fd_sc_hd__and2_1
XFILLER_30_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7360_ _7355_/A _7360_/B vssd1 vssd1 vccd1 vccd1 _7360_/X sky130_fd_sc_hd__and2b_1
X_4572_ _8582_/Q _8581_/Q _8584_/Q _8583_/Q vssd1 vssd1 vccd1 vccd1 _4573_/D sky130_fd_sc_hd__or4_1
X_7291_ _7307_/C _7291_/B vssd1 vssd1 vccd1 vccd1 _7377_/B sky130_fd_sc_hd__or2_1
X_6311_ _6311_/A _6311_/B vssd1 vssd1 vccd1 vccd1 _6312_/B sky130_fd_sc_hd__or2_1
XFILLER_6_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6242_ _6242_/A _6242_/B vssd1 vssd1 vccd1 vccd1 _6243_/B sky130_fd_sc_hd__xor2_2
XFILLER_97_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6173_ _5975_/A _6173_/B vssd1 vssd1 vccd1 vccd1 _6173_/X sky130_fd_sc_hd__and2b_1
XFILLER_84_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5124_ _5110_/B _5248_/C _5117_/X _5123_/X vssd1 vssd1 vccd1 vccd1 _5125_/A sky130_fd_sc_hd__o31a_1
X_5055_ _5172_/C _5055_/B _5055_/C vssd1 vssd1 vccd1 vccd1 _5055_/X sky130_fd_sc_hd__or3_1
XFILLER_72_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8796__74 vssd1 vssd1 vccd1 vccd1 _8796__74/HI _8905_/A sky130_fd_sc_hd__conb_1
XFILLER_25_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5957_ _6042_/B _5957_/B vssd1 vssd1 vccd1 vccd1 _5958_/A sky130_fd_sc_hd__or2_1
XFILLER_13_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4908_ _4908_/A vssd1 vssd1 vccd1 vccd1 _5011_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_8676_ input3/X _8676_/D vssd1 vssd1 vccd1 vccd1 _8676_/Q sky130_fd_sc_hd__dfxtp_1
X_7627_ _7627_/A _7627_/B vssd1 vssd1 vccd1 vccd1 _7673_/B sky130_fd_sc_hd__and2_1
X_5888_ _5990_/A _5888_/B vssd1 vssd1 vccd1 vccd1 _5916_/A sky130_fd_sc_hd__and2_1
X_4839_ _4839_/A _4839_/B vssd1 vssd1 vccd1 vccd1 _5094_/A sky130_fd_sc_hd__nor2_1
X_7558_ _8539_/B vssd1 vssd1 vccd1 vccd1 _8552_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_7489_ _7490_/A _7490_/B _7489_/C vssd1 vssd1 vccd1 vccd1 _7489_/X sky130_fd_sc_hd__or3_1
X_6509_ _5354_/B _6512_/A _6567_/A vssd1 vssd1 vccd1 vccd1 _6510_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6860_ _7202_/A vssd1 vssd1 vccd1 vccd1 _7151_/A sky130_fd_sc_hd__buf_2
X_6791_ _7176_/B _7176_/C vssd1 vssd1 vccd1 vccd1 _6919_/B sky130_fd_sc_hd__nand2_1
XFILLER_22_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5811_ _5812_/A _5812_/B vssd1 vssd1 vccd1 vccd1 _5887_/B sky130_fd_sc_hd__and2_1
X_5742_ _5742_/A _5742_/B vssd1 vssd1 vccd1 vccd1 _5920_/A sky130_fd_sc_hd__nor2_2
X_8530_ _8533_/A _7581_/X _8529_/Y vssd1 vssd1 vccd1 vccd1 _8719_/D sky130_fd_sc_hd__o21a_1
X_8461_ _8317_/A _7877_/A _7741_/Y vssd1 vssd1 vccd1 vccd1 _8462_/C sky130_fd_sc_hd__o21ai_1
X_5673_ _5763_/A vssd1 vssd1 vccd1 vccd1 _6193_/A sky130_fd_sc_hd__buf_2
X_8392_ _8392_/A _8392_/B vssd1 vssd1 vccd1 vccd1 _8400_/A sky130_fd_sc_hd__and2_1
X_7412_ _7413_/A _7412_/B _7412_/C vssd1 vssd1 vccd1 vccd1 _7449_/A sky130_fd_sc_hd__nand3_1
X_4624_ _8583_/Q _4623_/B _4607_/X vssd1 vssd1 vccd1 vccd1 _4625_/B sky130_fd_sc_hd__o21ai_1
X_7343_ _7343_/A _7343_/B vssd1 vssd1 vccd1 vccd1 _7345_/C sky130_fd_sc_hd__xnor2_1
X_4555_ _8621_/Q _4563_/B vssd1 vssd1 vccd1 vccd1 _4556_/A sky130_fd_sc_hd__and2_1
X_7274_ _7341_/A _7341_/B vssd1 vssd1 vccd1 vccd1 _7275_/A sky130_fd_sc_hd__nand2_1
X_4486_ _8609_/Q vssd1 vssd1 vccd1 vccd1 _7658_/B sky130_fd_sc_hd__clkbuf_4
X_6225_ _5540_/B _6227_/S _6007_/B _6007_/A vssd1 vssd1 vccd1 vccd1 _6228_/A sky130_fd_sc_hd__a22o_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6156_ _6303_/A _6303_/C vssd1 vssd1 vccd1 vccd1 _6304_/B sky130_fd_sc_hd__or2_1
XFILLER_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5107_ _5229_/D _5243_/B _5109_/B _5238_/A vssd1 vssd1 vccd1 vccd1 _5107_/X sky130_fd_sc_hd__or4_1
XFILLER_85_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6087_ _6087_/A _6087_/B vssd1 vssd1 vccd1 vccd1 _6088_/B sky130_fd_sc_hd__nand2_1
XFILLER_72_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5038_ _5166_/A _5166_/B _5057_/C _5091_/D vssd1 vssd1 vccd1 vccd1 _5038_/Y sky130_fd_sc_hd__nor4_1
XFILLER_26_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6989_ _6998_/A _6988_/B _6988_/C vssd1 vssd1 vccd1 vccd1 _6989_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8659_ input3/X _8659_/D vssd1 vssd1 vccd1 vccd1 _8659_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4340_ input1/X vssd1 vssd1 vccd1 vccd1 _4365_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_98_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6010_ _5895_/B _6224_/A _5898_/B _6009_/Y vssd1 vssd1 vccd1 vccd1 _6011_/B sky130_fd_sc_hd__a22o_1
XFILLER_67_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7961_ _8025_/B _7960_/C _7960_/A vssd1 vssd1 vccd1 vccd1 _7967_/B sky130_fd_sc_hd__a21o_1
X_8766__44 vssd1 vssd1 vccd1 vccd1 _8766__44/HI _8861_/A sky130_fd_sc_hd__conb_1
X_7892_ _7892_/A _7892_/B _7892_/C vssd1 vssd1 vccd1 vccd1 _7893_/B sky130_fd_sc_hd__or3_1
X_6912_ _7057_/B _6911_/C _6911_/A vssd1 vssd1 vccd1 vccd1 _6914_/B sky130_fd_sc_hd__a21o_1
X_6843_ _6979_/A _6843_/B vssd1 vssd1 vccd1 vccd1 _6848_/A sky130_fd_sc_hd__nor2_1
XFILLER_35_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6774_ _6751_/A _6842_/A _6847_/A vssd1 vssd1 vccd1 vccd1 _6954_/B sky130_fd_sc_hd__a21bo_1
XFILLER_22_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8513_ _7848_/A _8520_/B _7847_/A vssd1 vssd1 vccd1 vccd1 _8513_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5725_ _5881_/B _6005_/B vssd1 vssd1 vccd1 vccd1 _5809_/A sky130_fd_sc_hd__nor2_2
X_8444_ _8365_/A _8365_/B _8443_/X vssd1 vssd1 vccd1 vccd1 _8448_/A sky130_fd_sc_hd__a21o_1
X_5656_ _6042_/A _5962_/A vssd1 vssd1 vccd1 vccd1 _5974_/A sky130_fd_sc_hd__or2_2
X_4607_ _4607_/A vssd1 vssd1 vccd1 vccd1 _4607_/X sky130_fd_sc_hd__clkbuf_2
X_8375_ _8375_/A _8476_/A vssd1 vssd1 vccd1 vccd1 _8421_/A sky130_fd_sc_hd__xnor2_1
X_5587_ _6119_/A _5883_/A vssd1 vssd1 vccd1 vccd1 _5587_/Y sky130_fd_sc_hd__nor2_2
XFILLER_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7326_ _7326_/A _7326_/B vssd1 vssd1 vccd1 vccd1 _7373_/A sky130_fd_sc_hd__xor2_1
X_4538_ _4824_/B _4802_/B vssd1 vssd1 vccd1 vccd1 _4849_/B sky130_fd_sc_hd__nand2_2
X_7257_ _7268_/A _7268_/C _7268_/B vssd1 vssd1 vccd1 vccd1 _7260_/A sky130_fd_sc_hd__a21bo_1
X_4469_ _6560_/B vssd1 vssd1 vccd1 vccd1 _4705_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_77_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6208_ _6208_/A _6208_/B vssd1 vssd1 vccd1 vccd1 _6209_/B sky130_fd_sc_hd__nand2_1
X_7188_ _7188_/A _7173_/A vssd1 vssd1 vccd1 vccd1 _7188_/X sky130_fd_sc_hd__or2b_1
XFILLER_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6139_ _6140_/B _6140_/C _6140_/A vssd1 vssd1 vccd1 vccd1 _6303_/A sky130_fd_sc_hd__o21ai_2
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5510_ _5559_/B _5724_/B _5724_/C vssd1 vssd1 vccd1 vccd1 _5563_/A sky130_fd_sc_hd__and3_1
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6490_ _8703_/Q vssd1 vssd1 vccd1 vccd1 _7529_/A sky130_fd_sc_hd__clkbuf_2
X_5441_ _5441_/A _8646_/Q vssd1 vssd1 vccd1 vccd1 _5447_/B sky130_fd_sc_hd__or2_1
X_8160_ _8161_/A _8161_/B vssd1 vssd1 vccd1 vccd1 _8254_/B sky130_fd_sc_hd__and2_1
X_5372_ _8642_/Q _5373_/B vssd1 vssd1 vccd1 vccd1 _5374_/B sky130_fd_sc_hd__or2_1
X_7111_ _7031_/S _7107_/Y _7111_/S vssd1 vssd1 vccd1 vccd1 _7112_/B sky130_fd_sc_hd__mux2_1
X_8091_ _8263_/A _8263_/B vssd1 vssd1 vccd1 vccd1 _8499_/B sky130_fd_sc_hd__xnor2_1
X_7042_ _7042_/A _7042_/B vssd1 vssd1 vccd1 vccd1 _7078_/A sky130_fd_sc_hd__xnor2_1
XFILLER_86_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7944_ _7944_/A _7832_/B vssd1 vssd1 vccd1 vccd1 _8097_/A sky130_fd_sc_hd__or2b_2
XFILLER_55_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7875_ _7875_/A _6599_/B vssd1 vssd1 vccd1 vccd1 _7875_/X sky130_fd_sc_hd__or2b_1
X_6826_ _6771_/A _6771_/B _6825_/X vssd1 vssd1 vccd1 vccd1 _6851_/A sky130_fd_sc_hd__a21o_1
XFILLER_50_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6757_ _7184_/A _7184_/B vssd1 vssd1 vccd1 vccd1 _6757_/Y sky130_fd_sc_hd__nand2_1
XFILLER_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5708_ _5711_/B _5711_/C vssd1 vssd1 vccd1 vccd1 _5709_/C sky130_fd_sc_hd__nand2_1
X_6688_ _6642_/X _6643_/X _6657_/A vssd1 vssd1 vccd1 vccd1 _7047_/A sky130_fd_sc_hd__a21o_1
XFILLER_6_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8427_ _8427_/A _8427_/B vssd1 vssd1 vccd1 vccd1 _8493_/B sky130_fd_sc_hd__xor2_1
X_5639_ _5652_/A _5652_/B vssd1 vssd1 vccd1 vccd1 _5953_/B sky130_fd_sc_hd__xnor2_4
X_8358_ _8445_/A _8279_/B _8288_/B _8287_/B _8287_/A vssd1 vssd1 vccd1 vccd1 _8442_/A
+ sky130_fd_sc_hd__a32o_1
X_7309_ _7339_/A _7339_/B vssd1 vssd1 vccd1 vccd1 _7311_/B sky130_fd_sc_hd__xor2_1
XFILLER_2_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8289_ _8306_/A _8289_/B vssd1 vssd1 vccd1 vccd1 _8290_/B sky130_fd_sc_hd__xnor2_1
XFILLER_58_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5990_ _5990_/A _5990_/B vssd1 vssd1 vccd1 vccd1 _5991_/B sky130_fd_sc_hd__xor2_1
X_8736__14 vssd1 vssd1 vccd1 vccd1 _8736__14/HI _8831_/A sky130_fd_sc_hd__conb_1
X_4941_ _5238_/A _5153_/A _4941_/C _4940_/Y vssd1 vssd1 vccd1 vccd1 _4941_/X sky130_fd_sc_hd__or4b_1
X_7660_ _7660_/A _7660_/B vssd1 vssd1 vccd1 vccd1 _8305_/A sky130_fd_sc_hd__xnor2_4
X_4872_ _4872_/A _4872_/B _4872_/C vssd1 vssd1 vccd1 vccd1 _5026_/C sky130_fd_sc_hd__and3_1
X_6611_ _7193_/A _6806_/A vssd1 vssd1 vccd1 vccd1 _6751_/A sky130_fd_sc_hd__or2_2
XFILLER_20_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7591_ _8536_/A _7591_/B vssd1 vssd1 vccd1 vccd1 _7592_/A sky130_fd_sc_hd__and2_1
X_6542_ _6542_/A _6541_/X vssd1 vssd1 vccd1 vccd1 _6542_/X sky130_fd_sc_hd__or2b_1
XFILLER_9_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6473_ _8641_/Q _8640_/Q _6472_/X vssd1 vssd1 vccd1 vccd1 _6478_/C sky130_fd_sc_hd__or3b_1
X_8212_ _8212_/A _8212_/B _8212_/C vssd1 vssd1 vccd1 vccd1 _8213_/B sky130_fd_sc_hd__or3_1
X_5424_ _5425_/A _5425_/B vssd1 vssd1 vccd1 vccd1 _5424_/Y sky130_fd_sc_hd__nor2_1
X_8143_ _7786_/A _7786_/B _7644_/A _7644_/B _7908_/X vssd1 vssd1 vccd1 vccd1 _8305_/B
+ sky130_fd_sc_hd__a2111o_2
XFILLER_99_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5355_ _5355_/A vssd1 vssd1 vccd1 vccd1 _8636_/D sky130_fd_sc_hd__clkbuf_1
X_8074_ _8074_/A _8000_/B vssd1 vssd1 vccd1 vccd1 _8086_/A sky130_fd_sc_hd__or2b_1
X_5286_ _8617_/Q _5288_/B vssd1 vssd1 vccd1 vccd1 _5286_/X sky130_fd_sc_hd__or2_1
XINSDIODE2_6 _8522_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7025_ _7131_/A _7025_/B vssd1 vssd1 vccd1 vccd1 _7025_/X sky130_fd_sc_hd__and2_1
XFILLER_101_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7927_ _7927_/A _7927_/B vssd1 vssd1 vccd1 vccd1 _7928_/B sky130_fd_sc_hd__and2_1
XFILLER_55_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7858_ _7759_/A _7759_/B _7857_/X vssd1 vssd1 vccd1 vccd1 _7882_/A sky130_fd_sc_hd__a21o_1
X_6809_ _6737_/A _6737_/B _7194_/B _7092_/A vssd1 vssd1 vccd1 vccd1 _6947_/B sky130_fd_sc_hd__a211o_2
XFILLER_51_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7789_ _7789_/A _7789_/B vssd1 vssd1 vccd1 vccd1 _8302_/A sky130_fd_sc_hd__xor2_4
XFILLER_23_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8820__98 vssd1 vssd1 vccd1 vccd1 _8820__98/HI _8644_/D sky130_fd_sc_hd__conb_1
XFILLER_80_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5140_ _5253_/A _5137_/X _5139_/X _5070_/D _5149_/A vssd1 vssd1 vccd1 vccd1 _5140_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5071_ _5071_/A _5135_/D vssd1 vssd1 vccd1 vccd1 _5071_/X sky130_fd_sc_hd__or2_2
XFILLER_96_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8830_ _8830_/A _4338_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[9] sky130_fd_sc_hd__ebufn_8
X_5973_ _5971_/Y _5973_/B vssd1 vssd1 vccd1 vccd1 _5974_/B sky130_fd_sc_hd__and2b_1
XFILLER_25_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7712_ _7739_/A vssd1 vssd1 vccd1 vccd1 _7886_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4924_ _4923_/X _4990_/B vssd1 vssd1 vccd1 vccd1 _4928_/A sky130_fd_sc_hd__and2b_1
XFILLER_40_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8692_ input3/X _8692_/D vssd1 vssd1 vccd1 vccd1 _8692_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7643_ _7643_/A _7643_/B _7643_/C vssd1 vssd1 vccd1 vccd1 _7644_/B sky130_fd_sc_hd__and3_1
X_4855_ _5091_/A _5110_/B vssd1 vssd1 vccd1 vccd1 _5219_/C sky130_fd_sc_hd__or2_1
X_7574_ _8714_/Q vssd1 vssd1 vccd1 vccd1 _7574_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4786_ _5226_/A _4786_/B vssd1 vssd1 vccd1 vccd1 _5213_/B sky130_fd_sc_hd__or2_1
X_6525_ _6526_/A _6531_/B vssd1 vssd1 vccd1 vccd1 _6525_/Y sky130_fd_sc_hd__nor2_1
X_6456_ _6459_/C _6456_/B vssd1 vssd1 vccd1 vccd1 _8680_/D sky130_fd_sc_hd__nor2_1
X_5407_ _8557_/A _5419_/A vssd1 vssd1 vccd1 vccd1 _5412_/A sky130_fd_sc_hd__nor2_1
X_6387_ _8675_/Q _8674_/Q _8676_/Q vssd1 vssd1 vccd1 vccd1 _6387_/X sky130_fd_sc_hd__a21o_1
X_8126_ _8222_/A _8126_/B vssd1 vssd1 vccd1 vccd1 _8127_/B sky130_fd_sc_hd__xnor2_1
X_5338_ _8631_/Q _5336_/A _5325_/X vssd1 vssd1 vccd1 vccd1 _5339_/B sky130_fd_sc_hd__o21ai_1
X_8057_ _8057_/A _8280_/A _8057_/C _8057_/D vssd1 vssd1 vccd1 vccd1 _8172_/A sky130_fd_sc_hd__and4_1
XFILLER_87_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7008_ _7008_/A _7008_/B vssd1 vssd1 vccd1 vccd1 _7010_/C sky130_fd_sc_hd__xnor2_1
XFILLER_75_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5269_ _5269_/A _5269_/B _5269_/C vssd1 vssd1 vccd1 vccd1 _5269_/Y sky130_fd_sc_hd__nand3_1
XFILLER_47_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4640_ _4640_/A vssd1 vssd1 vccd1 vccd1 _8588_/D sky130_fd_sc_hd__clkbuf_1
X_6310_ _6310_/A _6310_/B vssd1 vssd1 vccd1 vccd1 _6310_/X sky130_fd_sc_hd__xor2_1
X_4571_ _6536_/B vssd1 vssd1 vccd1 vccd1 _4581_/A sky130_fd_sc_hd__clkbuf_4
X_7290_ _7231_/A _7376_/A _7230_/X vssd1 vssd1 vccd1 vccd1 _7291_/B sky130_fd_sc_hd__o21ba_1
X_6241_ _6241_/A _6246_/B vssd1 vssd1 vccd1 vccd1 _6242_/B sky130_fd_sc_hd__xnor2_2
X_6172_ _6027_/A _6027_/B _6171_/X vssd1 vssd1 vccd1 vccd1 _6242_/A sky130_fd_sc_hd__a21o_1
XFILLER_69_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5123_ _5176_/A _5231_/B _5123_/C _5256_/B vssd1 vssd1 vccd1 vccd1 _5123_/X sky130_fd_sc_hd__or4_1
XFILLER_69_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5054_ _5202_/A _5172_/B _5054_/C _5054_/D vssd1 vssd1 vccd1 vccd1 _5055_/C sky130_fd_sc_hd__or4_1
XFILLER_84_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5956_ _5956_/A _5956_/B vssd1 vssd1 vccd1 vccd1 _5986_/A sky130_fd_sc_hd__nor2_2
XFILLER_40_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4907_ _5231_/A _5092_/A _5215_/B _4907_/D vssd1 vssd1 vccd1 vccd1 _4907_/X sky130_fd_sc_hd__or4_1
X_8675_ input3/X _8675_/D vssd1 vssd1 vccd1 vccd1 _8675_/Q sky130_fd_sc_hd__dfxtp_1
X_5887_ _5887_/A _5887_/B _5887_/C vssd1 vssd1 vccd1 vccd1 _5888_/B sky130_fd_sc_hd__or3_1
X_7626_ _7627_/A _7627_/B vssd1 vssd1 vccd1 vccd1 _7673_/A sky130_fd_sc_hd__nor2_2
X_4838_ _4865_/B _4961_/A vssd1 vssd1 vccd1 vccd1 _5015_/A sky130_fd_sc_hd__nor2_1
XFILLER_21_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7557_ _8706_/Q vssd1 vssd1 vccd1 vccd1 _8539_/B sky130_fd_sc_hd__inv_2
X_4769_ _4769_/A vssd1 vssd1 vccd1 vccd1 _5263_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7488_ _7488_/A _7488_/B vssd1 vssd1 vccd1 vccd1 _7489_/C sky130_fd_sc_hd__nor2_1
X_6508_ _8688_/Q vssd1 vssd1 vccd1 vccd1 _6567_/A sky130_fd_sc_hd__inv_2
XFILLER_4_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6439_ _6441_/B _6441_/C _6419_/X vssd1 vssd1 vccd1 vccd1 _6439_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_20_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8109_ _8109_/A _8030_/A vssd1 vssd1 vccd1 vccd1 _8109_/X sky130_fd_sc_hd__or2b_1
XFILLER_102_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6790_ _6790_/A _6790_/B vssd1 vssd1 vccd1 vccd1 _6823_/B sky130_fd_sc_hd__nand2_1
X_5810_ _5810_/A _5879_/C vssd1 vssd1 vccd1 vccd1 _5812_/B sky130_fd_sc_hd__xnor2_1
X_5741_ _5600_/A _5599_/B _5740_/Y vssd1 vssd1 vccd1 vccd1 _5742_/B sky130_fd_sc_hd__o21a_1
X_8460_ _8460_/A _8460_/B vssd1 vssd1 vccd1 vccd1 _8464_/A sky130_fd_sc_hd__xnor2_1
X_7411_ _7409_/A _7409_/C _7409_/B vssd1 vssd1 vccd1 vccd1 _7412_/C sky130_fd_sc_hd__a21o_1
X_5672_ _6323_/C _5923_/B _5753_/A vssd1 vssd1 vccd1 vccd1 _5763_/A sky130_fd_sc_hd__mux2_2
X_8391_ _8343_/A _8343_/B _8342_/A vssd1 vssd1 vccd1 vccd1 _8453_/A sky130_fd_sc_hd__a21oi_1
X_4623_ _8583_/Q _4623_/B vssd1 vssd1 vccd1 vccd1 _4628_/C sky130_fd_sc_hd__and2_1
X_7342_ _7350_/A _7350_/B vssd1 vssd1 vccd1 vccd1 _7343_/B sky130_fd_sc_hd__xnor2_1
X_4554_ _4567_/B vssd1 vssd1 vccd1 vccd1 _4563_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_7273_ _7276_/A _7276_/B vssd1 vssd1 vccd1 vccd1 _7353_/A sky130_fd_sc_hd__xor2_1
XFILLER_103_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4485_ _4789_/A vssd1 vssd1 vccd1 vccd1 _4495_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6224_ _6224_/A vssd1 vssd1 vccd1 vccd1 _6227_/S sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_97_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6155_ _6303_/B _6303_/C vssd1 vssd1 vccd1 vccd1 _6316_/A sky130_fd_sc_hd__nor2_1
XFILLER_97_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5106_ _5087_/X _5103_/X _5014_/C _5104_/X _5105_/X vssd1 vssd1 vccd1 vccd1 _5106_/X
+ sky130_fd_sc_hd__o32a_1
X_6086_ _6087_/A _6087_/B vssd1 vssd1 vccd1 vccd1 _6094_/A sky130_fd_sc_hd__or2_1
X_5037_ _4823_/B _5026_/C _5241_/C vssd1 vssd1 vccd1 vccd1 _5166_/B sky130_fd_sc_hd__a21o_2
XFILLER_38_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6988_ _6998_/A _6988_/B _6988_/C vssd1 vssd1 vccd1 vccd1 _6988_/X sky130_fd_sc_hd__or3_2
XFILLER_13_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5939_ _5939_/A _5939_/B vssd1 vssd1 vccd1 vccd1 _5943_/B sky130_fd_sc_hd__xnor2_1
XFILLER_40_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8658_ input3/X _8658_/D vssd1 vssd1 vccd1 vccd1 _8658_/Q sky130_fd_sc_hd__dfxtp_2
X_7609_ _7604_/Y _7616_/B _7608_/X vssd1 vssd1 vccd1 vccd1 _7611_/C sky130_fd_sc_hd__a21oi_1
X_8589_ input3/X _8589_/D vssd1 vssd1 vccd1 vccd1 _8589_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7960_ _7960_/A _8025_/B _7960_/C vssd1 vssd1 vccd1 vccd1 _8023_/A sky130_fd_sc_hd__nand3_1
XFILLER_82_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7891_ _7892_/A _7892_/B _7892_/C vssd1 vssd1 vccd1 vccd1 _7980_/A sky130_fd_sc_hd__o21a_1
X_6911_ _6911_/A _7057_/B _6911_/C vssd1 vssd1 vccd1 vccd1 _6914_/A sky130_fd_sc_hd__nand3_1
XFILLER_54_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6842_ _6842_/A _6883_/B vssd1 vssd1 vccd1 vccd1 _6843_/B sky130_fd_sc_hd__and2_1
XFILLER_23_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8781__59 vssd1 vssd1 vccd1 vccd1 _8781__59/HI _8890_/A sky130_fd_sc_hd__conb_1
X_6773_ _6773_/A _7107_/A vssd1 vssd1 vccd1 vccd1 _6847_/A sky130_fd_sc_hd__nand2_2
XFILLER_62_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8512_ _8512_/A _8512_/B vssd1 vssd1 vccd1 vccd1 _8520_/B sky130_fd_sc_hd__nor2_1
X_5724_ _6009_/A _5724_/B _5724_/C vssd1 vssd1 vccd1 vccd1 _5726_/A sky130_fd_sc_hd__and3b_2
X_8443_ _8364_/A _8443_/B vssd1 vssd1 vccd1 vccd1 _8443_/X sky130_fd_sc_hd__and2b_1
X_5655_ _5957_/B vssd1 vssd1 vccd1 vccd1 _5962_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8374_ _7817_/X _8445_/A _8296_/B _8373_/Y vssd1 vssd1 vccd1 vccd1 _8476_/A sky130_fd_sc_hd__a31oi_2
X_4606_ _4610_/C _4606_/B vssd1 vssd1 vccd1 vccd1 _8577_/D sky130_fd_sc_hd__nor2_1
X_7325_ _7325_/A _7325_/B _7325_/C vssd1 vssd1 vccd1 vccd1 _7330_/A sky130_fd_sc_hd__nand3_1
X_5586_ _6005_/B vssd1 vssd1 vccd1 vccd1 _5883_/A sky130_fd_sc_hd__clkbuf_2
X_4537_ _4810_/A _4810_/B vssd1 vssd1 vccd1 vccd1 _4831_/C sky130_fd_sc_hd__nand2_1
XFILLER_104_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7256_ _7264_/A _7264_/B _7256_/C vssd1 vssd1 vccd1 vccd1 _7268_/B sky130_fd_sc_hd__nand3_1
X_4468_ _8597_/Q vssd1 vssd1 vccd1 vccd1 _6560_/B sky130_fd_sc_hd__buf_2
X_7187_ _7187_/A _7187_/B vssd1 vssd1 vccd1 vccd1 _7272_/B sky130_fd_sc_hd__xnor2_1
XFILLER_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6207_ _6207_/A _6207_/B _6207_/C vssd1 vssd1 vccd1 vccd1 _6208_/B sky130_fd_sc_hd__nand3_1
X_4399_ _4401_/A vssd1 vssd1 vccd1 vccd1 _4399_/Y sky130_fd_sc_hd__inv_2
X_6138_ _6138_/A _6149_/B vssd1 vssd1 vccd1 vccd1 _6140_/A sky130_fd_sc_hd__xnor2_1
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6069_ _6065_/A _6069_/B vssd1 vssd1 vccd1 vccd1 _6101_/A sky130_fd_sc_hd__and2b_1
XFILLER_85_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5440_ _5441_/A _8646_/Q vssd1 vssd1 vccd1 vccd1 _5442_/C sky130_fd_sc_hd__nand2_1
X_5371_ _5373_/B _5371_/B vssd1 vssd1 vccd1 vccd1 _8641_/D sky130_fd_sc_hd__nor2_1
X_7110_ _7195_/A _7110_/B vssd1 vssd1 vccd1 vccd1 _7111_/S sky130_fd_sc_hd__and2_1
X_8090_ _8090_/A _8090_/B vssd1 vssd1 vccd1 vccd1 _8263_/B sky130_fd_sc_hd__xor2_1
XFILLER_99_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7041_ _7041_/A vssd1 vssd1 vccd1 vccd1 _7042_/B sky130_fd_sc_hd__inv_2
XFILLER_86_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7943_ _8015_/A _7943_/B vssd1 vssd1 vccd1 vccd1 _8097_/B sky130_fd_sc_hd__or2_2
XFILLER_82_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7874_ _7885_/A _8115_/A vssd1 vssd1 vccd1 vccd1 _7964_/A sky130_fd_sc_hd__nor2_1
XFILLER_23_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6825_ _6785_/A _6825_/B vssd1 vssd1 vccd1 vccd1 _6825_/X sky130_fd_sc_hd__and2b_1
XFILLER_50_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6756_ _7184_/A _7184_/B vssd1 vssd1 vccd1 vccd1 _6756_/X sky130_fd_sc_hd__or2_1
XFILLER_23_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5707_ _6040_/A _6040_/B vssd1 vssd1 vccd1 vccd1 _5711_/C sky130_fd_sc_hd__or2_1
X_6687_ _6687_/A _6687_/B vssd1 vssd1 vccd1 vccd1 _6695_/A sky130_fd_sc_hd__xor2_1
X_8426_ _8439_/A _8426_/B vssd1 vssd1 vccd1 vccd1 _8427_/B sky130_fd_sc_hd__nor2_1
X_5638_ _5638_/A _5638_/B vssd1 vssd1 vccd1 vccd1 _5652_/B sky130_fd_sc_hd__nor2_2
X_8357_ _8312_/A _8312_/B _8313_/B _8313_/A vssd1 vssd1 vccd1 vccd1 _8477_/B sky130_fd_sc_hd__a2bb2o_1
X_5569_ _5569_/A _5569_/B _5568_/X vssd1 vssd1 vccd1 vccd1 _5576_/B sky130_fd_sc_hd__or3b_1
X_7308_ _7308_/A _7308_/B vssd1 vssd1 vccd1 vccd1 _7339_/B sky130_fd_sc_hd__nor2_1
XFILLER_2_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8288_ _8288_/A _8288_/B vssd1 vssd1 vccd1 vccd1 _8290_/A sky130_fd_sc_hd__xnor2_2
XFILLER_104_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7239_ _7239_/A _7239_/B vssd1 vssd1 vccd1 vccd1 _7241_/B sky130_fd_sc_hd__xor2_1
X_8726__4 vssd1 vssd1 vccd1 vccd1 _8726__4/HI _8821_/A sky130_fd_sc_hd__conb_1
XFILLER_58_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4940_ _5214_/D _5173_/B _5176_/C vssd1 vssd1 vccd1 vccd1 _4940_/Y sky130_fd_sc_hd__nor3_1
X_4871_ _4871_/A _4930_/B vssd1 vssd1 vccd1 vccd1 _5007_/A sky130_fd_sc_hd__nor2_1
XFILLER_32_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6610_ _6737_/A _6737_/B _6635_/A vssd1 vssd1 vccd1 vccd1 _6806_/A sky130_fd_sc_hd__a21o_2
X_7590_ _7589_/Y _7587_/A _8568_/A vssd1 vssd1 vccd1 vccd1 _7591_/B sky130_fd_sc_hd__mux2_1
X_8751__29 vssd1 vssd1 vccd1 vccd1 _8751__29/HI _8846_/A sky130_fd_sc_hd__conb_1
X_6541_ _6540_/A _6545_/A _6545_/B _6540_/D vssd1 vssd1 vccd1 vccd1 _6541_/X sky130_fd_sc_hd__a22o_1
X_6472_ _8639_/Q _8638_/Q _8643_/Q _8642_/Q vssd1 vssd1 vccd1 vccd1 _6472_/X sky130_fd_sc_hd__and4_1
X_8211_ _8212_/A _8212_/B _8212_/C vssd1 vssd1 vccd1 vccd1 _8312_/A sky130_fd_sc_hd__o21ai_2
X_5423_ _5414_/A _5421_/B _5415_/Y vssd1 vssd1 vccd1 vccd1 _5425_/B sky130_fd_sc_hd__a21oi_1
X_8142_ _8306_/B vssd1 vssd1 vccd1 vccd1 _8361_/A sky130_fd_sc_hd__clkbuf_2
X_5354_ _5360_/C _5354_/B _5354_/C vssd1 vssd1 vccd1 vccd1 _5355_/A sky130_fd_sc_hd__and3b_1
XFILLER_99_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8073_ _8073_/A _8101_/B vssd1 vssd1 vccd1 vccd1 _8088_/A sky130_fd_sc_hd__xnor2_1
X_5285_ _5285_/A vssd1 vssd1 vccd1 vccd1 _5285_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_59_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_7 _8534_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7024_ _7024_/A _7024_/B vssd1 vssd1 vccd1 vccd1 _7027_/A sky130_fd_sc_hd__xnor2_1
XFILLER_74_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7926_ _7927_/A _7927_/B vssd1 vssd1 vccd1 vccd1 _8018_/A sky130_fd_sc_hd__nor2_1
XFILLER_70_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7857_ _8209_/A _8218_/A _7857_/C vssd1 vssd1 vccd1 vccd1 _7857_/X sky130_fd_sc_hd__and3_1
XFILLER_23_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6808_ _7179_/A _7006_/A vssd1 vssd1 vccd1 vccd1 _6950_/A sky130_fd_sc_hd__nor2_2
XFILLER_51_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7788_ _7788_/A _8060_/B vssd1 vssd1 vccd1 vccd1 _7800_/A sky130_fd_sc_hd__nand2_1
XFILLER_11_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6739_ _7226_/A _7174_/B vssd1 vssd1 vccd1 vccd1 _7301_/A sky130_fd_sc_hd__nor2_4
XFILLER_11_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8409_ _8410_/A _8409_/B vssd1 vssd1 vccd1 vccd1 _8409_/X sky130_fd_sc_hd__or2_1
XFILLER_2_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5070_ _5214_/B _5214_/D _5149_/B _5070_/D vssd1 vssd1 vccd1 vccd1 _5070_/X sky130_fd_sc_hd__or4_1
XFILLER_56_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5972_ _5972_/A _5972_/B _5972_/C vssd1 vssd1 vccd1 vccd1 _5973_/B sky130_fd_sc_hd__nand3_1
XFILLER_18_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7711_ _7722_/A _7722_/B vssd1 vssd1 vccd1 vccd1 _7739_/A sky130_fd_sc_hd__xor2_1
X_4923_ _5110_/B _5193_/D vssd1 vssd1 vccd1 vccd1 _4923_/X sky130_fd_sc_hd__or2_1
X_8691_ input3/X _8691_/D vssd1 vssd1 vccd1 vccd1 _8691_/Q sky130_fd_sc_hd__dfxtp_1
X_7642_ _7643_/A _7643_/B _7643_/C vssd1 vssd1 vccd1 vccd1 _7644_/A sky130_fd_sc_hd__a21oi_1
X_4854_ _5042_/A _5240_/C vssd1 vssd1 vccd1 vccd1 _5110_/B sky130_fd_sc_hd__or2_2
XFILLER_33_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7573_ _7658_/A _7615_/B vssd1 vssd1 vccd1 vccd1 _7611_/A sky130_fd_sc_hd__nand2_1
X_4785_ _5226_/A _4786_/B vssd1 vssd1 vccd1 vccd1 _5213_/A sky130_fd_sc_hd__nand2_1
XFILLER_20_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6524_ _6520_/A _6511_/X _6513_/X _6523_/X vssd1 vssd1 vccd1 vccd1 _8690_/D sky130_fd_sc_hd__a22o_1
X_6455_ _8680_/Q _6454_/B _6409_/B vssd1 vssd1 vccd1 vccd1 _6456_/B sky130_fd_sc_hd__o21ai_1
X_5406_ _8591_/Q _5406_/B vssd1 vssd1 vccd1 vccd1 _5419_/A sky130_fd_sc_hd__and2_1
X_6386_ _6430_/A _8670_/Q _6385_/X _8672_/Q vssd1 vssd1 vccd1 vccd1 _6386_/X sky130_fd_sc_hd__a211o_1
X_8125_ _8125_/A _8326_/B vssd1 vssd1 vccd1 vccd1 _8222_/A sky130_fd_sc_hd__or2_2
X_5337_ _8631_/Q _8630_/Q _5337_/C vssd1 vssd1 vccd1 vccd1 _5342_/C sky130_fd_sc_hd__and3_1
XFILLER_0_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8056_ _8384_/A _8056_/B vssd1 vssd1 vccd1 vccd1 _8057_/D sky130_fd_sc_hd__or2_1
X_5268_ _4495_/A _4541_/B _4567_/B _5266_/Y _5267_/X vssd1 vssd1 vccd1 vccd1 _5269_/C
+ sky130_fd_sc_hd__o2111a_1
X_7007_ _7030_/B _6880_/A _7006_/X vssd1 vssd1 vccd1 vccd1 _7008_/B sky130_fd_sc_hd__a21oi_1
XFILLER_56_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5199_ _5199_/A _5199_/B vssd1 vssd1 vccd1 vccd1 _5199_/Y sky130_fd_sc_hd__nor2_1
XFILLER_71_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7909_ _7786_/A _7786_/B _7664_/A _7908_/X vssd1 vssd1 vccd1 vccd1 _7912_/B sky130_fd_sc_hd__a211o_1
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8889_ _8889_/A _4424_/Y vssd1 vssd1 vccd1 vccd1 io_out[36] sky130_fd_sc_hd__ebufn_8
XFILLER_24_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4570_ _6406_/A vssd1 vssd1 vccd1 vccd1 _6536_/B sky130_fd_sc_hd__clkbuf_4
X_6240_ _6240_/A _6240_/B vssd1 vssd1 vccd1 vccd1 _6246_/B sky130_fd_sc_hd__xor2_2
XFILLER_69_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6171_ _6026_/B _6171_/B vssd1 vssd1 vccd1 vccd1 _6171_/X sky130_fd_sc_hd__and2b_1
XFILLER_97_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5122_ _5122_/A _5122_/B vssd1 vssd1 vccd1 vccd1 _5256_/B sky130_fd_sc_hd__or2_1
XFILLER_97_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5053_ _5083_/A _5122_/A _5172_/B _5053_/D vssd1 vssd1 vccd1 vccd1 _5053_/X sky130_fd_sc_hd__or4_1
XFILLER_65_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5955_ _5953_/Y _6322_/A _5956_/B vssd1 vssd1 vccd1 vccd1 _5967_/A sky130_fd_sc_hd__o21ba_1
XFILLER_52_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4906_ _5030_/C _4895_/X _4901_/X _5151_/B _4905_/X vssd1 vssd1 vccd1 vccd1 _4907_/D
+ sky130_fd_sc_hd__o32a_1
X_8674_ input3/X _8674_/D vssd1 vssd1 vccd1 vccd1 _8674_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5886_ _5887_/A _5887_/B _5887_/C vssd1 vssd1 vccd1 vccd1 _5990_/A sky130_fd_sc_hd__o21ai_2
X_7625_ _7574_/X _7623_/Y _7624_/Y vssd1 vssd1 vccd1 vccd1 _8714_/D sky130_fd_sc_hd__a21oi_1
X_4837_ _4922_/A _4890_/A _5215_/B vssd1 vssd1 vccd1 vccd1 _5091_/A sky130_fd_sc_hd__or3_2
XFILLER_21_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7556_ _8539_/A _8531_/A _8546_/A vssd1 vssd1 vccd1 vccd1 _7556_/X sky130_fd_sc_hd__o21a_1
X_4768_ _6406_/A vssd1 vssd1 vccd1 vccd1 _7547_/A sky130_fd_sc_hd__clkbuf_2
X_7487_ _7490_/A _7490_/B _7488_/A vssd1 vssd1 vccd1 vccd1 _7487_/X sky130_fd_sc_hd__a21o_1
X_4699_ _6556_/B _4699_/B vssd1 vssd1 vccd1 vccd1 _4994_/B sky130_fd_sc_hd__nor2_1
X_6507_ _6507_/A _7545_/B vssd1 vssd1 vccd1 vccd1 _6512_/A sky130_fd_sc_hd__nor2_1
XFILLER_20_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6438_ _6441_/C _6438_/B vssd1 vssd1 vccd1 vccd1 _8674_/D sky130_fd_sc_hd__nor2_1
XFILLER_88_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8108_ _8041_/A _8041_/B _8107_/Y vssd1 vssd1 vccd1 vccd1 _8133_/A sky130_fd_sc_hd__o21a_1
XFILLER_88_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6369_ _6367_/A _6376_/S vssd1 vssd1 vccd1 vccd1 _6373_/A sky130_fd_sc_hd__and2b_1
XFILLER_88_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8039_ _8039_/A _8039_/B vssd1 vssd1 vccd1 vccd1 _8040_/B sky130_fd_sc_hd__nor2_1
XFILLER_48_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8787__65 vssd1 vssd1 vccd1 vccd1 _8787__65/HI _8896_/A sky130_fd_sc_hd__conb_1
XFILLER_16_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5740_ _5740_/A _5740_/B vssd1 vssd1 vccd1 vccd1 _5740_/Y sky130_fd_sc_hd__nand2_1
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7410_ _7443_/A _6880_/A _7289_/B _7301_/A vssd1 vssd1 vccd1 vccd1 _7412_/B sky130_fd_sc_hd__a22o_1
X_5671_ _5671_/A _5957_/B vssd1 vssd1 vccd1 vccd1 _5753_/A sky130_fd_sc_hd__or2_2
X_8390_ _8390_/A _8390_/B vssd1 vssd1 vccd1 vccd1 _8419_/A sky130_fd_sc_hd__xnor2_1
X_4622_ _4622_/A vssd1 vssd1 vccd1 vccd1 _8582_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4553_ _4553_/A vssd1 vssd1 vccd1 vccd1 _8874_/A sky130_fd_sc_hd__clkbuf_1
X_7341_ _7341_/A _7341_/B vssd1 vssd1 vccd1 vccd1 _7350_/B sky130_fd_sc_hd__xnor2_1
X_7272_ _7272_/A _7272_/B vssd1 vssd1 vccd1 vccd1 _7276_/B sky130_fd_sc_hd__xnor2_1
X_4484_ _7631_/B vssd1 vssd1 vccd1 vccd1 _4789_/A sky130_fd_sc_hd__clkbuf_2
X_6223_ _6019_/A _6019_/B _6018_/A vssd1 vssd1 vccd1 vccd1 _6234_/A sky130_fd_sc_hd__a21bo_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6154_ _6163_/A _6164_/C vssd1 vssd1 vccd1 vccd1 _6303_/C sky130_fd_sc_hd__or2b_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5105_ _5105_/A vssd1 vssd1 vccd1 vccd1 _5105_/X sky130_fd_sc_hd__buf_2
X_6085_ _6085_/A _6085_/B vssd1 vssd1 vccd1 vccd1 _6134_/A sky130_fd_sc_hd__xnor2_1
XFILLER_85_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5036_ _5185_/A vssd1 vssd1 vccd1 vccd1 _5040_/A sky130_fd_sc_hd__inv_2
XFILLER_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6987_ _6987_/A _6987_/B vssd1 vssd1 vccd1 vccd1 _6988_/C sky130_fd_sc_hd__xnor2_1
XFILLER_80_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5938_ _5938_/A _5938_/B vssd1 vssd1 vccd1 vccd1 _5939_/B sky130_fd_sc_hd__xnor2_1
XFILLER_25_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5869_ _5983_/B _5870_/B vssd1 vssd1 vccd1 vccd1 _5869_/Y sky130_fd_sc_hd__nand2_1
X_8657_ input3/X _8657_/D vssd1 vssd1 vccd1 vccd1 _8657_/Q sky130_fd_sc_hd__dfxtp_1
X_7608_ _7604_/Y _7616_/B _7603_/B vssd1 vssd1 vccd1 vccd1 _7608_/X sky130_fd_sc_hd__o21a_1
X_8588_ input3/X _8588_/D vssd1 vssd1 vccd1 vccd1 _8588_/Q sky130_fd_sc_hd__dfxtp_1
X_7539_ _7539_/A _7539_/B vssd1 vssd1 vccd1 vccd1 _7540_/B sky130_fd_sc_hd__xnor2_1
XFILLER_31_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7890_ _8044_/A _7890_/B vssd1 vssd1 vccd1 vccd1 _7892_/C sky130_fd_sc_hd__and2_1
X_6910_ _7057_/A _6909_/C _7135_/A vssd1 vssd1 vccd1 vccd1 _6911_/C sky130_fd_sc_hd__a21o_1
XFILLER_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6841_ _6842_/A _6883_/B vssd1 vssd1 vccd1 vccd1 _6979_/A sky130_fd_sc_hd__nor2_1
XFILLER_35_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6772_ _6772_/A vssd1 vssd1 vccd1 vccd1 _7107_/A sky130_fd_sc_hd__buf_2
X_8511_ _8508_/A _8508_/B _7842_/C vssd1 vssd1 vccd1 vccd1 _8512_/B sky130_fd_sc_hd__a21oi_1
X_5723_ _6214_/A _5574_/B _5731_/A _5582_/B vssd1 vssd1 vccd1 vccd1 _5792_/A sky130_fd_sc_hd__a22o_1
X_8442_ _8442_/A _8442_/B vssd1 vssd1 vccd1 vccd1 _8442_/Y sky130_fd_sc_hd__nand2_1
X_5654_ _5616_/B _5629_/B _5759_/A vssd1 vssd1 vccd1 vccd1 _5957_/B sky130_fd_sc_hd__a21bo_1
X_8373_ _8294_/A _8294_/B _8295_/A vssd1 vssd1 vccd1 vccd1 _8373_/Y sky130_fd_sc_hd__a21oi_1
X_4605_ _8577_/Q _4603_/A _4595_/X vssd1 vssd1 vccd1 vccd1 _4606_/B sky130_fd_sc_hd__o21ai_1
XFILLER_30_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7324_ _7323_/B _7323_/C _7323_/A vssd1 vssd1 vccd1 vccd1 _7325_/C sky130_fd_sc_hd__a21o_1
X_5585_ _6323_/B _6005_/B vssd1 vssd1 vccd1 vccd1 _5795_/A sky130_fd_sc_hd__or2_1
X_4536_ _8602_/Q vssd1 vssd1 vccd1 vccd1 _4810_/B sky130_fd_sc_hd__inv_2
X_7255_ _7264_/A _7264_/B _7256_/C vssd1 vssd1 vccd1 vccd1 _7268_/C sky130_fd_sc_hd__a21o_1
X_4467_ _6605_/B vssd1 vssd1 vccd1 vccd1 _5226_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_4398_ _4401_/A vssd1 vssd1 vccd1 vccd1 _4398_/Y sky130_fd_sc_hd__inv_2
X_7186_ _7262_/B _7186_/B vssd1 vssd1 vccd1 vccd1 _7187_/B sky130_fd_sc_hd__xnor2_1
XFILLER_89_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6206_ _6207_/A _6207_/B _6207_/C vssd1 vssd1 vccd1 vccd1 _6208_/A sky130_fd_sc_hd__a21o_1
X_6137_ _6153_/A _6137_/B vssd1 vssd1 vccd1 vccd1 _6149_/B sky130_fd_sc_hd__and2b_1
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6068_ _6070_/B _6070_/A vssd1 vssd1 vccd1 vccd1 _6103_/A sky130_fd_sc_hd__and2b_1
X_8757__35 vssd1 vssd1 vccd1 vccd1 _8757__35/HI _8852_/A sky130_fd_sc_hd__conb_1
X_5019_ _5241_/C vssd1 vssd1 vccd1 vccd1 _5239_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_26_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8709_ input3/X _8709_/D vssd1 vssd1 vccd1 vccd1 _8709_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_9_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5370_ _8641_/Q _5369_/B _5357_/X vssd1 vssd1 vccd1 vccd1 _5371_/B sky130_fd_sc_hd__o21ai_1
XFILLER_99_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7040_ _7038_/Y _6961_/B _7039_/Y vssd1 vssd1 vccd1 vccd1 _7041_/A sky130_fd_sc_hd__a21oi_1
XFILLER_86_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7942_ _7942_/A _7942_/B _7942_/C vssd1 vssd1 vccd1 vccd1 _7943_/B sky130_fd_sc_hd__and3_1
XFILLER_70_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7873_ _7954_/B vssd1 vssd1 vccd1 vccd1 _8115_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6824_ _6824_/A _6824_/B vssd1 vssd1 vccd1 vccd1 _6895_/A sky130_fd_sc_hd__nand2_1
XFILLER_50_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6755_ _7180_/A _7313_/A _7266_/A vssd1 vssd1 vccd1 vccd1 _7184_/B sky130_fd_sc_hd__a21oi_1
X_5706_ _5706_/A _5706_/B vssd1 vssd1 vccd1 vccd1 _6040_/B sky130_fd_sc_hd__xnor2_1
X_8425_ _8425_/A _8425_/B _8425_/C vssd1 vssd1 vccd1 vccd1 _8426_/B sky130_fd_sc_hd__nor3_1
X_6686_ _6614_/X _6642_/X _6643_/X _6798_/A _7238_/A vssd1 vssd1 vccd1 vccd1 _6689_/A
+ sky130_fd_sc_hd__a311oi_1
X_5637_ _5680_/A vssd1 vssd1 vccd1 vccd1 _5638_/A sky130_fd_sc_hd__inv_2
X_8356_ _8347_/A _8347_/B _8355_/X vssd1 vssd1 vccd1 vccd1 _8482_/A sky130_fd_sc_hd__a21o_1
X_5568_ _5603_/A _5568_/B vssd1 vssd1 vccd1 vccd1 _5568_/X sky130_fd_sc_hd__and2b_1
X_7307_ _7307_/A _7307_/B _7307_/C vssd1 vssd1 vccd1 vccd1 _7308_/B sky130_fd_sc_hd__nor3_1
X_8287_ _8287_/A _8287_/B vssd1 vssd1 vccd1 vccd1 _8288_/B sky130_fd_sc_hd__xor2_2
X_4519_ _6599_/B _7753_/A vssd1 vssd1 vccd1 vccd1 _4732_/A sky130_fd_sc_hd__nand2_1
XFILLER_104_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7238_ _7238_/A _7297_/B _7299_/B vssd1 vssd1 vccd1 vccd1 _7241_/A sky130_fd_sc_hd__or3_1
X_5499_ _5499_/A vssd1 vssd1 vccd1 vccd1 _5559_/B sky130_fd_sc_hd__buf_2
XFILLER_104_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7169_ _7169_/A _7169_/B _7169_/C vssd1 vssd1 vccd1 vccd1 _7262_/B sky130_fd_sc_hd__nand3_4
XFILLER_85_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4870_ _4898_/B vssd1 vssd1 vccd1 vccd1 _4930_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_60_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6540_ _6540_/A _6545_/A _6545_/B _6540_/D vssd1 vssd1 vccd1 vccd1 _6542_/A sky130_fd_sc_hd__and4_1
X_6471_ _8631_/Q _8630_/Q _6471_/C _8634_/Q vssd1 vssd1 vccd1 vccd1 _6478_/B sky130_fd_sc_hd__nand4_1
X_8210_ _8462_/B _8475_/A _8381_/A vssd1 vssd1 vccd1 vccd1 _8212_/C sky130_fd_sc_hd__o21a_1
X_5422_ _5422_/A _5422_/B vssd1 vssd1 vccd1 vccd1 _5425_/A sky130_fd_sc_hd__or2_1
X_8141_ _8141_/A _8152_/A vssd1 vssd1 vccd1 vccd1 _8306_/B sky130_fd_sc_hd__nand2_1
X_5353_ _6471_/C _8634_/Q _5346_/B _8636_/Q vssd1 vssd1 vccd1 vccd1 _5354_/C sky130_fd_sc_hd__a31o_1
X_8072_ _8072_/A _8072_/B vssd1 vssd1 vccd1 vccd1 _8101_/B sky130_fd_sc_hd__xor2_1
X_5284_ _8715_/Q _5271_/X _5282_/X _5283_/X vssd1 vssd1 vccd1 vccd1 _8616_/D sky130_fd_sc_hd__o211a_1
XFILLER_87_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7023_ _7023_/A _7118_/B vssd1 vssd1 vccd1 vccd1 _7024_/B sky130_fd_sc_hd__xor2_1
XINSDIODE2_8 _6617_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7925_ _7801_/A _7801_/B _7924_/Y vssd1 vssd1 vccd1 vccd1 _7927_/B sky130_fd_sc_hd__a21oi_1
X_7856_ _7856_/A vssd1 vssd1 vccd1 vccd1 _8218_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_70_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6807_ _6807_/A vssd1 vssd1 vccd1 vccd1 _7006_/A sky130_fd_sc_hd__buf_2
X_7787_ _7911_/B vssd1 vssd1 vccd1 vccd1 _8060_/B sky130_fd_sc_hd__buf_2
X_4999_ _4952_/A _4987_/X _4993_/X _5190_/A _5190_/C vssd1 vssd1 vccd1 vccd1 _4999_/X
+ sky130_fd_sc_hd__a311o_1
X_6738_ _6863_/A vssd1 vssd1 vccd1 vccd1 _7174_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_7_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6669_ _7238_/A _6798_/B _7237_/C _7177_/A _7245_/B vssd1 vssd1 vccd1 vccd1 _6670_/A
+ sky130_fd_sc_hd__o32ai_2
X_8408_ _8408_/A _8408_/B vssd1 vssd1 vccd1 vccd1 _8412_/A sky130_fd_sc_hd__xor2_1
X_8339_ _8404_/A _8404_/B vssd1 vssd1 vccd1 vccd1 _8341_/C sky130_fd_sc_hd__xnor2_1
XFILLER_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8811__89 vssd1 vssd1 vccd1 vccd1 _8811__89/HI _8920_/A sky130_fd_sc_hd__conb_1
X_5971_ _5972_/A _5972_/B _5972_/C vssd1 vssd1 vccd1 vccd1 _5971_/Y sky130_fd_sc_hd__a21oi_1
X_7710_ _7746_/A _7823_/A vssd1 vssd1 vccd1 vccd1 _7885_/A sky130_fd_sc_hd__nand2_2
X_4922_ _4922_/A _4937_/C vssd1 vssd1 vccd1 vccd1 _5193_/D sky130_fd_sc_hd__or2_2
XFILLER_18_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8690_ input3/X _8690_/D vssd1 vssd1 vccd1 vccd1 _8690_/Q sky130_fd_sc_hd__dfxtp_1
X_7641_ _7639_/X _7641_/B vssd1 vssd1 vccd1 vccd1 _7643_/C sky130_fd_sc_hd__and2b_1
XFILLER_33_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4853_ _5041_/A _5041_/B _5017_/A vssd1 vssd1 vccd1 vccd1 _5240_/C sky130_fd_sc_hd__o21ai_2
X_7572_ _8712_/Q vssd1 vssd1 vccd1 vccd1 _7658_/A sky130_fd_sc_hd__inv_2
X_4784_ _4784_/A _4784_/B vssd1 vssd1 vccd1 vccd1 _8611_/D sky130_fd_sc_hd__nor2_1
X_6523_ _6523_/A _6523_/B vssd1 vssd1 vccd1 vccd1 _6523_/X sky130_fd_sc_hd__xor2_1
X_6454_ _8680_/Q _6454_/B vssd1 vssd1 vccd1 vccd1 _6459_/C sky130_fd_sc_hd__and2_1
X_5405_ _6507_/A vssd1 vssd1 vccd1 vccd1 _8557_/A sky130_fd_sc_hd__buf_2
X_6385_ _8667_/Q _8668_/Q _8671_/Q _6397_/D vssd1 vssd1 vccd1 vccd1 _6385_/X sky130_fd_sc_hd__o211a_1
X_8124_ _8317_/A _8462_/A vssd1 vssd1 vccd1 vccd1 _8127_/A sky130_fd_sc_hd__nor2_1
X_5336_ _5336_/A _5336_/B vssd1 vssd1 vccd1 vccd1 _8630_/D sky130_fd_sc_hd__nor2_1
X_8055_ _8168_/C _8055_/B vssd1 vssd1 vccd1 vccd1 _8057_/C sky130_fd_sc_hd__and2_1
X_5267_ _4782_/A _4781_/A _4769_/A _4535_/C _4775_/A vssd1 vssd1 vccd1 vccd1 _5267_/X
+ sky130_fd_sc_hd__o221a_1
X_7006_ _7006_/A _7031_/S _7065_/B vssd1 vssd1 vccd1 vccd1 _7006_/X sky130_fd_sc_hd__and3_1
XFILLER_68_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5198_ _4885_/X _5151_/A _5137_/B _5176_/D _5166_/D vssd1 vssd1 vccd1 vccd1 _5199_/B
+ sky130_fd_sc_hd__o41a_1
XFILLER_18_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7908_ _7574_/X _7908_/B vssd1 vssd1 vccd1 vccd1 _7908_/X sky130_fd_sc_hd__and2b_1
X_8888_ _8888_/A _4426_/Y vssd1 vssd1 vccd1 vccd1 io_out[35] sky130_fd_sc_hd__ebufn_8
XFILLER_24_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7839_ _7839_/A _7839_/B vssd1 vssd1 vccd1 vccd1 _8206_/A sky130_fd_sc_hd__nor2_1
XFILLER_70_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6170_ _6170_/A _6028_/B vssd1 vssd1 vccd1 vccd1 _6244_/A sky130_fd_sc_hd__or2b_1
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5121_ _5116_/B _5193_/A _5118_/X _5120_/X vssd1 vssd1 vccd1 vccd1 _5123_/C sky130_fd_sc_hd__o31a_1
XFILLER_69_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5052_ _5166_/A vssd1 vssd1 vccd1 vccd1 _5214_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_37_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5954_ _5954_/A _5954_/B _5954_/C vssd1 vssd1 vccd1 vccd1 _6322_/A sky130_fd_sc_hd__and3_2
X_4905_ _4989_/A _5098_/B _4976_/B _5074_/B vssd1 vssd1 vccd1 vccd1 _4905_/X sky130_fd_sc_hd__or4_1
X_8673_ input3/X _8673_/D vssd1 vssd1 vccd1 vccd1 _8673_/Q sky130_fd_sc_hd__dfxtp_1
X_5885_ _5993_/A _6263_/A _6259_/A vssd1 vssd1 vccd1 vccd1 _5887_/C sky130_fd_sc_hd__mux2_1
X_7624_ _7574_/X _7623_/Y _4581_/A vssd1 vssd1 vccd1 vccd1 _7624_/Y sky130_fd_sc_hd__o21ai_1
X_4836_ _4861_/A _4836_/B vssd1 vssd1 vccd1 vccd1 _5215_/B sky130_fd_sc_hd__nor2_2
XFILLER_21_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7555_ _8722_/Q vssd1 vssd1 vccd1 vccd1 _8546_/A sky130_fd_sc_hd__clkbuf_2
X_6506_ _6500_/X _6505_/Y _5273_/X vssd1 vssd1 vccd1 vccd1 _8687_/D sky130_fd_sc_hd__o21ai_1
X_4767_ _4767_/A vssd1 vssd1 vccd1 vccd1 _8607_/D sky130_fd_sc_hd__clkbuf_1
X_7486_ _7486_/A _7486_/B _7486_/C vssd1 vssd1 vccd1 vccd1 _7492_/C sky130_fd_sc_hd__or3_1
X_4698_ _6556_/B _7708_/B _8594_/Q vssd1 vssd1 vccd1 vccd1 _4994_/A sky130_fd_sc_hd__and3_1
X_6437_ _8674_/Q _6435_/A _6409_/B vssd1 vssd1 vccd1 vccd1 _6438_/B sky130_fd_sc_hd__o21ai_1
XFILLER_20_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6368_ _5413_/A _6366_/Y _6376_/S _5412_/X _8662_/Q vssd1 vssd1 vccd1 vccd1 _8662_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_96_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8107_ _8107_/A _8107_/B vssd1 vssd1 vccd1 vccd1 _8107_/Y sky130_fd_sc_hd__nand2_1
X_5319_ _8626_/Q _8625_/Q _8624_/Q vssd1 vssd1 vccd1 vccd1 _5324_/B sky130_fd_sc_hd__and3_1
XFILLER_88_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6299_ _6299_/A _6299_/B vssd1 vssd1 vccd1 vccd1 _6341_/A sky130_fd_sc_hd__xnor2_4
XFILLER_102_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8038_ _8109_/A _8038_/B vssd1 vssd1 vccd1 vccd1 _8039_/B sky130_fd_sc_hd__and2_1
XFILLER_75_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5670_ _5754_/A _6110_/B vssd1 vssd1 vccd1 vccd1 _5674_/A sky130_fd_sc_hd__nand2_2
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4621_ _4623_/B _4639_/B _4621_/C vssd1 vssd1 vccd1 vccd1 _4622_/A sky130_fd_sc_hd__and3b_1
X_7340_ _7323_/A _7323_/C _7323_/B vssd1 vssd1 vccd1 vccd1 _7350_/A sky130_fd_sc_hd__a21boi_2
X_4552_ _8620_/Q _4552_/B vssd1 vssd1 vccd1 vccd1 _4553_/A sky130_fd_sc_hd__and2_1
X_7271_ _7336_/B _7336_/C _7336_/D _7270_/X vssd1 vssd1 vccd1 vccd1 _7276_/A sky130_fd_sc_hd__o31a_1
X_4483_ _8606_/Q vssd1 vssd1 vccd1 vccd1 _7631_/B sky130_fd_sc_hd__clkbuf_4
X_6222_ _6222_/A _6222_/B vssd1 vssd1 vccd1 vccd1 _6266_/A sky130_fd_sc_hd__xnor2_2
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6153_ _6153_/A _6153_/B _6151_/Y vssd1 vssd1 vccd1 vccd1 _6164_/C sky130_fd_sc_hd__or3b_1
XFILLER_97_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5104_ _5110_/B _5104_/B _5256_/A _5202_/B vssd1 vssd1 vccd1 vccd1 _5104_/X sky130_fd_sc_hd__or4_1
X_6084_ _6085_/A _6085_/B vssd1 vssd1 vccd1 vccd1 _6084_/X sky130_fd_sc_hd__or2_1
XFILLER_85_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5035_ _5149_/A _5193_/D _5022_/X _5034_/X _4953_/X vssd1 vssd1 vccd1 vccd1 _5060_/C
+ sky130_fd_sc_hd__o311a_1
XFILLER_53_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6986_ _6996_/B _6986_/B vssd1 vssd1 vccd1 vccd1 _6987_/B sky130_fd_sc_hd__xnor2_1
X_8725_ input3/X _8725_/D vssd1 vssd1 vccd1 vccd1 _8725_/Q sky130_fd_sc_hd__dfxtp_1
X_5937_ _5937_/A _5937_/B vssd1 vssd1 vccd1 vccd1 _5938_/B sky130_fd_sc_hd__nand2_1
X_8656_ input3/X _8656_/D vssd1 vssd1 vccd1 vccd1 _8656_/Q sky130_fd_sc_hd__dfxtp_1
X_7607_ _7658_/A _7616_/B vssd1 vssd1 vccd1 vccd1 _7611_/B sky130_fd_sc_hd__or2_1
X_5868_ _5844_/A _5844_/B _5867_/Y vssd1 vssd1 vccd1 vccd1 _5946_/A sky130_fd_sc_hd__a21oi_1
X_4819_ _4872_/C _4872_/A vssd1 vssd1 vccd1 vccd1 _4820_/B sky130_fd_sc_hd__and2b_1
X_8587_ input3/X _8587_/D vssd1 vssd1 vccd1 vccd1 _8587_/Q sky130_fd_sc_hd__dfxtp_1
X_5799_ _5801_/C _6034_/B vssd1 vssd1 vccd1 vccd1 _6213_/B sky130_fd_sc_hd__nand2_1
X_7538_ _7543_/B _7538_/B vssd1 vssd1 vccd1 vccd1 _7539_/B sky130_fd_sc_hd__nand2_1
X_7469_ _7469_/A _7469_/B vssd1 vssd1 vccd1 vccd1 _7492_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6840_ _6863_/A _6864_/A vssd1 vssd1 vccd1 vccd1 _6883_/B sky130_fd_sc_hd__or2_2
X_6771_ _6771_/A _6771_/B vssd1 vssd1 vccd1 vccd1 _6785_/A sky130_fd_sc_hd__xnor2_1
XFILLER_50_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8510_ _8527_/A _8527_/B _8520_/A vssd1 vssd1 vccd1 vccd1 _8510_/X sky130_fd_sc_hd__and3_1
X_5722_ _5720_/X _5590_/B _5721_/X vssd1 vssd1 vccd1 vccd1 _5789_/A sky130_fd_sc_hd__a21o_1
XFILLER_50_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8441_ _8441_/A _8366_/B vssd1 vssd1 vccd1 vccd1 _8441_/X sky130_fd_sc_hd__or2b_1
X_5653_ _5666_/A _5961_/A vssd1 vssd1 vccd1 vccd1 _5704_/A sky130_fd_sc_hd__nand2_1
X_8372_ _8477_/B _8372_/B vssd1 vssd1 vccd1 vccd1 _8375_/A sky130_fd_sc_hd__xnor2_1
X_4604_ _8576_/Q _8577_/Q _4604_/C vssd1 vssd1 vccd1 vccd1 _4610_/C sky130_fd_sc_hd__and3_1
X_5584_ _5584_/A _5584_/B vssd1 vssd1 vccd1 vccd1 _6323_/B sky130_fd_sc_hd__and2_1
X_7323_ _7323_/A _7323_/B _7323_/C vssd1 vssd1 vccd1 vccd1 _7325_/B sky130_fd_sc_hd__nand3_1
XFILLER_7_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4535_ _4775_/A _4769_/A _4535_/C vssd1 vssd1 vccd1 vccd1 _4541_/B sky130_fd_sc_hd__nand3_1
XFILLER_104_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7254_ _7254_/A _7254_/B vssd1 vssd1 vccd1 vccd1 _7256_/C sky130_fd_sc_hd__xor2_1
X_4466_ _7699_/B vssd1 vssd1 vccd1 vccd1 _6605_/B sky130_fd_sc_hd__clkbuf_2
X_4397_ _4401_/A vssd1 vssd1 vccd1 vccd1 _4397_/Y sky130_fd_sc_hd__inv_2
X_7185_ _7185_/A _7185_/B vssd1 vssd1 vccd1 vccd1 _7186_/B sky130_fd_sc_hd__xnor2_1
X_6205_ _6205_/A _6269_/B vssd1 vssd1 vccd1 vccd1 _6207_/C sky130_fd_sc_hd__xnor2_1
X_6136_ _6135_/A _6135_/C _6135_/B vssd1 vssd1 vccd1 vccd1 _6137_/B sky130_fd_sc_hd__o21ai_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6067_ _6097_/A _6097_/B _6066_/X vssd1 vssd1 vccd1 vccd1 _6070_/A sky130_fd_sc_hd__a21o_1
XFILLER_85_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5018_ _5118_/B _5182_/C _4916_/B _5191_/A _5143_/B vssd1 vssd1 vccd1 vccd1 _5018_/X
+ sky130_fd_sc_hd__o41a_1
XFILLER_45_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6969_ _7151_/A _6891_/B _6968_/X vssd1 vssd1 vccd1 vccd1 _6987_/A sky130_fd_sc_hd__a21o_1
XFILLER_53_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8708_ input3/X _8708_/D vssd1 vssd1 vccd1 vccd1 _8708_/Q sky130_fd_sc_hd__dfxtp_1
X_8639_ input3/X _8639_/D vssd1 vssd1 vccd1 vccd1 _8639_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7941_ _7942_/A _7942_/B _7942_/C vssd1 vssd1 vccd1 vccd1 _8015_/A sky130_fd_sc_hd__a21oi_1
XFILLER_67_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7872_ _7766_/A _7871_/X _7766_/C _7751_/A vssd1 vssd1 vccd1 vccd1 _7954_/B sky130_fd_sc_hd__a31o_1
XFILLER_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6823_ _6823_/A _6823_/B _6823_/C vssd1 vssd1 vccd1 vccd1 _6824_/B sky130_fd_sc_hd__nand3_1
XFILLER_90_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6754_ _7239_/A _6842_/A vssd1 vssd1 vccd1 vccd1 _7266_/A sky130_fd_sc_hd__nor2_2
XFILLER_11_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6685_ _6685_/A vssd1 vssd1 vccd1 vccd1 _6719_/A sky130_fd_sc_hd__buf_2
XFILLER_50_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5705_ _6063_/B _5705_/B vssd1 vssd1 vccd1 vccd1 _5706_/B sky130_fd_sc_hd__nor2_1
X_8424_ _8425_/A _8425_/B _8425_/C vssd1 vssd1 vccd1 vccd1 _8439_/A sky130_fd_sc_hd__o21a_1
XFILLER_12_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5636_ _5657_/A _5657_/B _5622_/X vssd1 vssd1 vccd1 vccd1 _5652_/A sky130_fd_sc_hd__a21o_2
XFILLER_31_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8355_ _8346_/A _8355_/B vssd1 vssd1 vccd1 vccd1 _8355_/X sky130_fd_sc_hd__and2b_1
X_5567_ _5567_/A _5567_/B _5567_/C vssd1 vssd1 vccd1 vccd1 _5568_/B sky130_fd_sc_hd__or3_1
X_7306_ _7306_/A _7306_/B vssd1 vssd1 vccd1 vccd1 _7339_/A sky130_fd_sc_hd__xnor2_1
X_8286_ _8301_/B _8360_/B _8286_/C vssd1 vssd1 vccd1 vccd1 _8287_/B sky130_fd_sc_hd__and3_1
X_4518_ _7908_/B _5617_/A _4518_/C _4660_/B vssd1 vssd1 vccd1 vccd1 _4520_/B sky130_fd_sc_hd__or4_1
X_5498_ _5584_/A _5584_/B vssd1 vssd1 vccd1 vccd1 _5499_/A sky130_fd_sc_hd__nand2_1
X_4449_ _4450_/A vssd1 vssd1 vccd1 vccd1 _4449_/Y sky130_fd_sc_hd__inv_2
X_7237_ _7245_/A _7237_/B _7237_/C vssd1 vssd1 vccd1 vccd1 _7299_/B sky130_fd_sc_hd__or3_2
X_8817__95 vssd1 vssd1 vccd1 vccd1 _8817__95/HI _8926_/A sky130_fd_sc_hd__conb_1
X_7168_ _7168_/A _7168_/B vssd1 vssd1 vccd1 vccd1 _7169_/C sky130_fd_sc_hd__xnor2_2
XFILLER_100_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7099_ _7099_/A _7099_/B vssd1 vssd1 vccd1 vccd1 _7100_/B sky130_fd_sc_hd__xnor2_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6119_ _6119_/A _6119_/B vssd1 vssd1 vccd1 vccd1 _6121_/B sky130_fd_sc_hd__xnor2_1
XFILLER_100_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6470_ _8705_/Q vssd1 vssd1 vccd1 vccd1 _7545_/A sky130_fd_sc_hd__inv_2
X_5421_ _5421_/A _5421_/B vssd1 vssd1 vccd1 vccd1 _5422_/B sky130_fd_sc_hd__nor2_1
X_8140_ _8140_/A _8140_/B vssd1 vssd1 vccd1 vccd1 _8161_/A sky130_fd_sc_hd__nor2_1
X_5352_ _8636_/Q _6471_/C _5352_/C vssd1 vssd1 vccd1 vccd1 _5360_/C sky130_fd_sc_hd__and3_1
X_8071_ _8071_/A _8071_/B vssd1 vssd1 vccd1 vccd1 _8072_/B sky130_fd_sc_hd__xnor2_1
XFILLER_99_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7022_ _7133_/A _7022_/B vssd1 vssd1 vccd1 vccd1 _7118_/B sky130_fd_sc_hd__nand2_1
XFILLER_59_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5283_ _5296_/A vssd1 vssd1 vccd1 vccd1 _5283_/X sky130_fd_sc_hd__clkbuf_2
XINSDIODE2_9 _7783_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7924_ _7924_/A _7924_/B vssd1 vssd1 vccd1 vccd1 _7924_/Y sky130_fd_sc_hd__nor2_1
XFILLER_36_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7855_ _8125_/A vssd1 vssd1 vccd1 vccd1 _7856_/A sky130_fd_sc_hd__inv_2
XFILLER_63_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6806_ _6806_/A _6806_/B vssd1 vssd1 vccd1 vccd1 _6807_/A sky130_fd_sc_hd__or2_1
XFILLER_23_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7786_ _7786_/A _7786_/B vssd1 vssd1 vccd1 vccd1 _7911_/B sky130_fd_sc_hd__xor2_1
XFILLER_51_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4998_ _5139_/A vssd1 vssd1 vccd1 vccd1 _5190_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_6737_ _6737_/A _6737_/B vssd1 vssd1 vccd1 vccd1 _6863_/A sky130_fd_sc_hd__xnor2_2
XFILLER_23_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6668_ _7175_/B vssd1 vssd1 vccd1 vccd1 _7245_/B sky130_fd_sc_hd__clkbuf_2
X_8407_ _7964_/X _8406_/Y _8407_/S vssd1 vssd1 vccd1 vccd1 _8408_/B sky130_fd_sc_hd__mux2_1
X_6599_ _7545_/A _6599_/B vssd1 vssd1 vccd1 vccd1 _6600_/B sky130_fd_sc_hd__nor2_1
X_5619_ _6617_/A _8650_/Q vssd1 vssd1 vccd1 vccd1 _5679_/A sky130_fd_sc_hd__or2b_1
X_8338_ _8415_/A _8338_/B vssd1 vssd1 vccd1 vccd1 _8404_/B sky130_fd_sc_hd__and2_1
XFILLER_2_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8269_ _8269_/A _8269_/B vssd1 vssd1 vccd1 vccd1 _8269_/Y sky130_fd_sc_hd__nor2_1
XFILLER_59_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5970_ _6190_/B _5970_/B vssd1 vssd1 vccd1 vccd1 _5972_/C sky130_fd_sc_hd__xor2_1
XFILLER_37_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4921_ _4930_/A _4836_/B _4834_/X vssd1 vssd1 vccd1 vccd1 _4937_/C sky130_fd_sc_hd__o21ai_4
X_7640_ _8608_/Q _8711_/Q vssd1 vssd1 vccd1 vccd1 _7641_/B sky130_fd_sc_hd__or2b_1
X_4852_ _5227_/B _5026_/B _5046_/A vssd1 vssd1 vccd1 vccd1 _5017_/A sky130_fd_sc_hd__a21oi_2
X_7571_ _7594_/A _7571_/B vssd1 vssd1 vccd1 vccd1 _7571_/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4783_ _4782_/A _5275_/B _4782_/Y _4739_/B vssd1 vssd1 vccd1 vccd1 _4784_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_9_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6522_ _6514_/A _6526_/B _6515_/Y vssd1 vssd1 vccd1 vccd1 _6523_/B sky130_fd_sc_hd__a21o_1
X_6453_ _6453_/A vssd1 vssd1 vccd1 vccd1 _8679_/D sky130_fd_sc_hd__clkbuf_1
X_5404_ _5402_/C _5398_/Y _5403_/Y _5296_/X vssd1 vssd1 vccd1 vccd1 _8646_/D sky130_fd_sc_hd__o211a_1
X_8123_ _8326_/B vssd1 vssd1 vccd1 vccd1 _8462_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6384_ _8669_/Q vssd1 vssd1 vccd1 vccd1 _6397_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_87_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5335_ _8630_/Q _5337_/C _5325_/X vssd1 vssd1 vccd1 vccd1 _5336_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8054_ _8054_/A _8054_/B vssd1 vssd1 vccd1 vccd1 _8055_/B sky130_fd_sc_hd__nand2_1
X_5266_ _5127_/B _5261_/C _4723_/X _5265_/X vssd1 vssd1 vccd1 vccd1 _5266_/Y sky130_fd_sc_hd__o31ai_1
X_7005_ _7236_/B _6954_/B _6847_/A vssd1 vssd1 vccd1 vccd1 _7008_/A sky130_fd_sc_hd__o21ai_1
XFILLER_68_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5197_ _5040_/A _4673_/A _5138_/Y _5196_/X _4727_/A vssd1 vssd1 vccd1 vccd1 _5197_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_28_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7907_ _8051_/A _8384_/A vssd1 vssd1 vccd1 vccd1 _7920_/A sky130_fd_sc_hd__nand2_1
XFILLER_70_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8887_ _8887_/A _4458_/Y vssd1 vssd1 vccd1 vccd1 io_out[34] sky130_fd_sc_hd__ebufn_8
XFILLER_70_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7838_ _8209_/A _8134_/A vssd1 vssd1 vccd1 vccd1 _7839_/B sky130_fd_sc_hd__nor2_1
XFILLER_24_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7769_ _7769_/A vssd1 vssd1 vccd1 vccd1 _8327_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_11_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5120_ _5120_/A _5231_/C _5120_/C _5120_/D vssd1 vssd1 vccd1 vccd1 _5120_/X sky130_fd_sc_hd__or4_1
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5051_ _5143_/A vssd1 vssd1 vccd1 vccd1 _5229_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_38_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5953_ _6123_/A _5953_/B vssd1 vssd1 vccd1 vccd1 _5953_/Y sky130_fd_sc_hd__nor2_1
X_4904_ _5159_/B _5152_/B vssd1 vssd1 vccd1 vccd1 _4976_/B sky130_fd_sc_hd__or2_1
X_5884_ _5997_/A _6323_/B _5907_/B vssd1 vssd1 vccd1 vccd1 _6263_/A sky130_fd_sc_hd__mux2_2
X_8672_ input3/X _8672_/D vssd1 vssd1 vccd1 vccd1 _8672_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7623_ _8564_/A _7623_/B vssd1 vssd1 vccd1 vccd1 _7623_/Y sky130_fd_sc_hd__nor2_1
XFILLER_60_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4835_ _4836_/B _4898_/A _4834_/X vssd1 vssd1 vccd1 vccd1 _4890_/A sky130_fd_sc_hd__o21ai_1
X_7554_ _8720_/Q vssd1 vssd1 vccd1 vccd1 _8531_/A sky130_fd_sc_hd__clkbuf_2
X_4766_ _4775_/C _7503_/A _4766_/C vssd1 vssd1 vccd1 vccd1 _4767_/A sky130_fd_sc_hd__and3b_1
X_6505_ _6505_/A _6505_/B vssd1 vssd1 vccd1 vccd1 _6505_/Y sky130_fd_sc_hd__nor2_1
X_7485_ _7485_/A _7485_/B vssd1 vssd1 vccd1 vccd1 _7486_/C sky130_fd_sc_hd__xor2_1
XFILLER_20_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4697_ _4970_/A _4697_/B vssd1 vssd1 vccd1 vccd1 _4697_/Y sky130_fd_sc_hd__nor2_1
X_6436_ _8674_/Q _8673_/Q _6436_/C vssd1 vssd1 vccd1 vccd1 _6441_/C sky130_fd_sc_hd__and3_1
X_6367_ _6367_/A _6367_/B _6367_/C vssd1 vssd1 vccd1 vccd1 _6376_/S sky130_fd_sc_hd__or3_1
X_8106_ _8047_/A _8047_/B _8105_/X vssd1 vssd1 vccd1 vccd1 _8191_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5318_ _5318_/A vssd1 vssd1 vccd1 vccd1 _8625_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6298_ _6298_/A _6298_/B vssd1 vssd1 vccd1 vccd1 _6299_/B sky130_fd_sc_hd__xnor2_4
X_8037_ _8109_/A _8038_/B vssd1 vssd1 vccd1 vccd1 _8039_/A sky130_fd_sc_hd__nor2_1
X_5249_ _5110_/D _5241_/X _5246_/X _5248_/X vssd1 vssd1 vccd1 vccd1 _5249_/X sky130_fd_sc_hd__o31a_1
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8778__56 vssd1 vssd1 vccd1 vccd1 _8778__56/HI _8887_/A sky130_fd_sc_hd__conb_1
XFILLER_74_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4620_ _8580_/Q _8581_/Q _4614_/B _8582_/Q vssd1 vssd1 vccd1 vccd1 _4621_/C sky130_fd_sc_hd__a31o_1
X_4551_ _4551_/A vssd1 vssd1 vccd1 vccd1 _8869_/A sky130_fd_sc_hd__clkbuf_2
X_7270_ _7270_/A _7313_/B _7334_/C _7334_/D vssd1 vssd1 vccd1 vccd1 _7270_/X sky130_fd_sc_hd__or4bb_1
X_4482_ _4850_/A vssd1 vssd1 vccd1 vccd1 _4745_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6221_ _5997_/A _5997_/B _6220_/X vssd1 vssd1 vccd1 vccd1 _6222_/B sky130_fd_sc_hd__a21oi_2
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6152_ _6153_/A _6153_/B _6151_/Y vssd1 vssd1 vccd1 vccd1 _6163_/A sky130_fd_sc_hd__o21ba_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5103_ _5122_/B _5103_/B vssd1 vssd1 vccd1 vccd1 _5103_/X sky130_fd_sc_hd__or2_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6083_ _6323_/A _6213_/A _6083_/C vssd1 vssd1 vccd1 vccd1 _6085_/B sky130_fd_sc_hd__or3_1
XFILLER_85_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5034_ _5159_/A _5034_/B vssd1 vssd1 vccd1 vccd1 _5034_/X sky130_fd_sc_hd__or2_1
X_6985_ _7205_/A _6985_/B vssd1 vssd1 vccd1 vccd1 _6986_/B sky130_fd_sc_hd__xnor2_1
XFILLER_53_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8724_ input3/X _8724_/D vssd1 vssd1 vccd1 vccd1 _8724_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5936_ _5936_/A _5936_/B vssd1 vssd1 vccd1 vccd1 _5938_/A sky130_fd_sc_hd__nor2_1
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8792__70 vssd1 vssd1 vccd1 vccd1 _8792__70/HI _8901_/A sky130_fd_sc_hd__conb_1
X_8655_ input3/X _8655_/D vssd1 vssd1 vccd1 vccd1 _8655_/Q sky130_fd_sc_hd__dfxtp_1
X_7606_ _7583_/X _7602_/X _7603_/Y _7605_/Y vssd1 vssd1 vccd1 vccd1 _8711_/D sky130_fd_sc_hd__o31a_1
XFILLER_21_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5867_ _5867_/A _5867_/B vssd1 vssd1 vccd1 vccd1 _5867_/Y sky130_fd_sc_hd__nor2_1
X_4818_ _4859_/A _4860_/A vssd1 vssd1 vccd1 vccd1 _4922_/A sky130_fd_sc_hd__nor2_1
XFILLER_21_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8586_ input3/X _8586_/D vssd1 vssd1 vccd1 vccd1 _8586_/Q sky130_fd_sc_hd__dfxtp_1
X_5798_ _5883_/A vssd1 vssd1 vccd1 vccd1 _6215_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7537_ _7537_/A _7537_/B vssd1 vssd1 vccd1 vccd1 _7538_/B sky130_fd_sc_hd__or2_1
XFILLER_5_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4749_ _6536_/B vssd1 vssd1 vccd1 vccd1 _8536_/A sky130_fd_sc_hd__clkbuf_2
X_7468_ _7490_/A _7490_/B _7465_/Y _7466_/X _7467_/X vssd1 vssd1 vccd1 vccd1 _7469_/B
+ sky130_fd_sc_hd__a32o_2
X_6419_ _6419_/A vssd1 vssd1 vccd1 vccd1 _6419_/X sky130_fd_sc_hd__clkbuf_2
X_7399_ _7399_/A _7399_/B vssd1 vssd1 vccd1 vccd1 _7402_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6770_ _6768_/X _7266_/A _6769_/X vssd1 vssd1 vccd1 vccd1 _6771_/B sky130_fd_sc_hd__o21ba_1
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5721_ _5721_/A _5721_/B vssd1 vssd1 vccd1 vccd1 _5721_/X sky130_fd_sc_hd__and2_1
XFILLER_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8440_ _8370_/A _8370_/B _8371_/B _8371_/A vssd1 vssd1 vccd1 vccd1 _8451_/A sky130_fd_sc_hd__o22a_1
X_5652_ _5652_/A _5652_/B vssd1 vssd1 vccd1 vccd1 _5961_/A sky130_fd_sc_hd__xor2_2
XFILLER_30_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8371_ _8371_/A _8371_/B vssd1 vssd1 vccd1 vccd1 _8372_/B sky130_fd_sc_hd__xnor2_1
X_5583_ _5721_/A _5721_/B vssd1 vssd1 vccd1 vccd1 _5590_/A sky130_fd_sc_hd__xnor2_1
X_4603_ _4603_/A _4603_/B vssd1 vssd1 vccd1 vccd1 _8576_/D sky130_fd_sc_hd__nor2_1
X_7322_ _7326_/A _7326_/B _7321_/C vssd1 vssd1 vccd1 vccd1 _7323_/C sky130_fd_sc_hd__a21o_1
X_4534_ _4723_/A _7753_/A _4534_/C _4662_/B vssd1 vssd1 vccd1 vccd1 _4542_/C sky130_fd_sc_hd__or4b_1
XFILLER_7_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7253_ _7250_/X _7318_/B _7252_/Y vssd1 vssd1 vccd1 vccd1 _7264_/B sky130_fd_sc_hd__a21bo_2
X_4465_ _8598_/Q vssd1 vssd1 vccd1 vccd1 _7699_/B sky130_fd_sc_hd__clkbuf_2
X_4396_ _4396_/A vssd1 vssd1 vccd1 vccd1 _4401_/A sky130_fd_sc_hd__buf_4
X_7184_ _7184_/A _7184_/B vssd1 vssd1 vccd1 vccd1 _7185_/B sky130_fd_sc_hd__xnor2_1
X_6204_ _6204_/A _6204_/B vssd1 vssd1 vccd1 vccd1 _6269_/B sky130_fd_sc_hd__or2_1
X_6135_ _6135_/A _6135_/B _6135_/C vssd1 vssd1 vccd1 vccd1 _6153_/A sky130_fd_sc_hd__nor3_1
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6066_ _6062_/A _6066_/B vssd1 vssd1 vccd1 vccd1 _6066_/X sky130_fd_sc_hd__and2b_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5017_ _5017_/A _5017_/B vssd1 vssd1 vccd1 vccd1 _5191_/A sky130_fd_sc_hd__nand2_1
XFILLER_66_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6968_ _6890_/B _6968_/B vssd1 vssd1 vccd1 vccd1 _6968_/X sky130_fd_sc_hd__and2b_1
X_8707_ input3/X _8707_/D vssd1 vssd1 vccd1 vccd1 _8707_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6899_ _6899_/A _7131_/A vssd1 vssd1 vccd1 vccd1 _6911_/A sky130_fd_sc_hd__and2_1
X_5919_ _5946_/A _5946_/B vssd1 vssd1 vccd1 vccd1 _5939_/A sky130_fd_sc_hd__xor2_1
X_8638_ input3/X _8638_/D vssd1 vssd1 vccd1 vccd1 _8638_/Q sky130_fd_sc_hd__dfxtp_1
X_8569_ _7875_/A _8568_/Y _4581_/A vssd1 vssd1 vccd1 vccd1 _8569_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_5_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8748__26 vssd1 vssd1 vccd1 vccd1 _8748__26/HI _8843_/A sky130_fd_sc_hd__conb_1
XFILLER_29_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7940_ _7940_/A _7940_/B vssd1 vssd1 vccd1 vccd1 _7942_/C sky130_fd_sc_hd__or2_1
XFILLER_82_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7871_ _7871_/A _8725_/Q vssd1 vssd1 vccd1 vccd1 _7871_/X sky130_fd_sc_hd__or2b_1
X_6822_ _6823_/A _6823_/B _6823_/C vssd1 vssd1 vccd1 vccd1 _6824_/A sky130_fd_sc_hd__a21o_1
XFILLER_63_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8762__40 vssd1 vssd1 vccd1 vccd1 _8762__40/HI _8857_/A sky130_fd_sc_hd__conb_1
X_6753_ _6947_/A _6753_/B vssd1 vssd1 vccd1 vccd1 _7313_/A sky130_fd_sc_hd__xor2_4
XFILLER_50_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6684_ _7418_/A _6919_/A vssd1 vssd1 vccd1 vccd1 _6685_/A sky130_fd_sc_hd__nor2_1
X_5704_ _5704_/A _5704_/B vssd1 vssd1 vccd1 vccd1 _5705_/B sky130_fd_sc_hd__and2_1
X_8423_ _8423_/A _8423_/B vssd1 vssd1 vccd1 vccd1 _8425_/C sky130_fd_sc_hd__xor2_1
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5635_ _5826_/A _5666_/A vssd1 vssd1 vccd1 vccd1 _5959_/A sky130_fd_sc_hd__nand2_1
X_8354_ _8298_/A _8298_/B _8353_/X vssd1 vssd1 vccd1 vccd1 _8423_/A sky130_fd_sc_hd__a21oi_1
X_5566_ _5567_/A _5567_/B _5567_/C vssd1 vssd1 vccd1 vccd1 _5603_/A sky130_fd_sc_hd__o21a_1
X_7305_ _7305_/A _7320_/A vssd1 vssd1 vccd1 vccd1 _7306_/B sky130_fd_sc_hd__xnor2_1
X_8285_ _8284_/C _8360_/A _7671_/A vssd1 vssd1 vccd1 vccd1 _8286_/C sky130_fd_sc_hd__a21o_1
X_4517_ _7658_/B _4769_/A _4535_/C _4789_/A vssd1 vssd1 vccd1 vccd1 _4660_/B sky130_fd_sc_hd__or4_1
X_5497_ _6343_/S _8595_/Q vssd1 vssd1 vccd1 vccd1 _5584_/B sky130_fd_sc_hd__nand2_1
XFILLER_104_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4448_ _4450_/A vssd1 vssd1 vccd1 vccd1 _4448_/Y sky130_fd_sc_hd__inv_2
X_7236_ _7236_/A _7236_/B vssd1 vssd1 vccd1 vccd1 _7320_/A sky130_fd_sc_hd__nor2_2
XFILLER_86_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7167_ _6697_/X _7167_/B vssd1 vssd1 vccd1 vccd1 _7168_/B sky130_fd_sc_hd__and2b_1
XFILLER_58_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4379_ _4383_/A vssd1 vssd1 vccd1 vccd1 _4379_/Y sky130_fd_sc_hd__inv_2
X_7098_ _7107_/A _7131_/A vssd1 vssd1 vccd1 vccd1 _7099_/B sky130_fd_sc_hd__xnor2_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6118_ _6323_/A _6083_/C _5800_/X vssd1 vssd1 vccd1 vccd1 _6119_/B sky130_fd_sc_hd__o21a_1
XFILLER_100_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6049_ _6049_/A _6049_/B vssd1 vssd1 vccd1 vccd1 _6050_/B sky130_fd_sc_hd__xnor2_1
XFILLER_37_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5420_ _5421_/A _5421_/B vssd1 vssd1 vccd1 vccd1 _5422_/A sky130_fd_sc_hd__and2_1
X_5351_ _6471_/C _5352_/C _5350_/Y vssd1 vssd1 vccd1 vccd1 _8635_/D sky130_fd_sc_hd__a21oi_1
XFILLER_99_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8070_ _8070_/A _8070_/B vssd1 vssd1 vccd1 vccd1 _8071_/B sky130_fd_sc_hd__nand2_1
X_5282_ _8616_/Q _5288_/B vssd1 vssd1 vccd1 vccd1 _5282_/X sky130_fd_sc_hd__or2_1
XFILLER_99_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7021_ _7065_/B _7179_/A vssd1 vssd1 vccd1 vccd1 _7022_/B sky130_fd_sc_hd__or2b_1
XFILLER_101_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7923_ _7923_/A _7923_/B vssd1 vssd1 vccd1 vccd1 _7927_/A sky130_fd_sc_hd__xnor2_1
XFILLER_82_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7854_ _7772_/A _7772_/B _7853_/X vssd1 vssd1 vccd1 vccd1 _7949_/A sky130_fd_sc_hd__a21o_1
XFILLER_36_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6805_ _6805_/A _6951_/A vssd1 vssd1 vccd1 vccd1 _6896_/A sky130_fd_sc_hd__or2b_1
X_7785_ _7679_/A _7676_/X _7679_/B _7677_/A vssd1 vssd1 vccd1 vccd1 _7786_/B sky130_fd_sc_hd__a31o_2
X_6736_ _6978_/A vssd1 vssd1 vccd1 vccd1 _7030_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_51_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4997_ _5135_/D vssd1 vssd1 vccd1 vccd1 _5139_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_23_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6667_ _6674_/A _6674_/B vssd1 vssd1 vccd1 vccd1 _7175_/B sky130_fd_sc_hd__xor2_2
X_8406_ _8406_/A _8406_/B vssd1 vssd1 vccd1 vccd1 _8406_/Y sky130_fd_sc_hd__nor2_1
X_6598_ _7545_/A _7871_/A vssd1 vssd1 vccd1 vccd1 _6635_/A sky130_fd_sc_hd__and2_1
X_5618_ _7658_/B _8651_/Q vssd1 vssd1 vccd1 vccd1 _5642_/A sky130_fd_sc_hd__or2b_1
X_8337_ _8410_/A _8337_/B _8409_/B vssd1 vssd1 vccd1 vccd1 _8338_/B sky130_fd_sc_hd__nand3_1
XFILLER_3_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5549_ _5549_/A _6599_/B vssd1 vssd1 vccd1 vccd1 _5549_/Y sky130_fd_sc_hd__nand2_1
XFILLER_2_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8268_ _8262_/A _8497_/B _8262_/B vssd1 vssd1 vccd1 vccd1 _8492_/C sky130_fd_sc_hd__o21ai_1
X_8199_ _8385_/A _8199_/B vssd1 vssd1 vccd1 vccd1 _8200_/B sky130_fd_sc_hd__and2_1
X_7219_ _7219_/A _7254_/A vssd1 vssd1 vccd1 vccd1 _7220_/B sky130_fd_sc_hd__xnor2_1
XFILLER_86_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4920_ _5071_/A _5238_/A _5098_/D _5137_/B vssd1 vssd1 vccd1 vccd1 _4920_/X sky130_fd_sc_hd__or4_1
XFILLER_33_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4851_ _4859_/A _5010_/B vssd1 vssd1 vccd1 vccd1 _5046_/A sky130_fd_sc_hd__nor2_2
XFILLER_60_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8732__10 vssd1 vssd1 vccd1 vccd1 _8732__10/HI _8827_/A sky130_fd_sc_hd__conb_1
X_7570_ _7587_/A _8708_/Q _7604_/A vssd1 vssd1 vccd1 vccd1 _7571_/B sky130_fd_sc_hd__a21oi_1
X_4782_ _4782_/A _4782_/B vssd1 vssd1 vccd1 vccd1 _4782_/Y sky130_fd_sc_hd__xnor2_1
X_6521_ _6521_/A _6521_/B vssd1 vssd1 vccd1 vccd1 _6523_/A sky130_fd_sc_hd__nor2_1
X_6452_ _6454_/B _6468_/B _6452_/C vssd1 vssd1 vccd1 vccd1 _6453_/A sky130_fd_sc_hd__and3b_1
X_5403_ _5433_/B _5403_/B vssd1 vssd1 vccd1 vccd1 _5403_/Y sky130_fd_sc_hd__nand2_1
X_8122_ _8205_/A _8205_/B vssd1 vssd1 vccd1 vccd1 _8128_/A sky130_fd_sc_hd__nand2_1
X_6383_ _8671_/Q vssd1 vssd1 vccd1 vccd1 _6430_/A sky130_fd_sc_hd__clkbuf_1
X_5334_ _8630_/Q _5337_/C vssd1 vssd1 vccd1 vccd1 _5336_/A sky130_fd_sc_hd__and2_1
XFILLER_102_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8053_ _8054_/A _8054_/B vssd1 vssd1 vccd1 vccd1 _8168_/C sky130_fd_sc_hd__or2_1
X_5265_ _5265_/A _6777_/B _5265_/C _4723_/A vssd1 vssd1 vccd1 vccd1 _5265_/X sky130_fd_sc_hd__or4b_1
XFILLER_87_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7004_ _7004_/A _7010_/A _7004_/C vssd1 vssd1 vccd1 vccd1 _7010_/B sky130_fd_sc_hd__nand3_1
X_5196_ _5144_/B _5203_/A _5192_/Y _5075_/Y _5195_/Y vssd1 vssd1 vccd1 vccd1 _5196_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_18_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8886_ _8886_/A _4407_/Y vssd1 vssd1 vccd1 vccd1 io_out[33] sky130_fd_sc_hd__ebufn_8
X_7906_ _8301_/A vssd1 vssd1 vccd1 vccd1 _8384_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_36_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7837_ _7864_/A vssd1 vssd1 vccd1 vccd1 _8209_/A sky130_fd_sc_hd__buf_2
XFILLER_24_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7768_ _7957_/C _7957_/D vssd1 vssd1 vccd1 vccd1 _7769_/A sky130_fd_sc_hd__nor2_1
X_6719_ _6719_/A _6814_/A vssd1 vssd1 vccd1 vccd1 _6900_/A sky130_fd_sc_hd__xnor2_2
X_7699_ _8722_/Q _7699_/B vssd1 vssd1 vccd1 vccd1 _7701_/A sky130_fd_sc_hd__and2b_1
XFILLER_50_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5050_ _5219_/B _5040_/X _5049_/X vssd1 vssd1 vccd1 vccd1 _5050_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5952_ _6323_/D _5923_/B _5926_/B _5951_/Y vssd1 vssd1 vccd1 vccd1 _6190_/B sky130_fd_sc_hd__a31o_1
XFILLER_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4903_ _4903_/A _4930_/B vssd1 vssd1 vccd1 vccd1 _5152_/B sky130_fd_sc_hd__nor2_1
XFILLER_18_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5883_ _5883_/A _6143_/B vssd1 vssd1 vccd1 vccd1 _5907_/B sky130_fd_sc_hd__nor2_1
X_8671_ input3/X _8671_/D vssd1 vssd1 vccd1 vccd1 _8671_/Q sky130_fd_sc_hd__dfxtp_1
X_7622_ _7621_/X _7617_/A _7622_/S vssd1 vssd1 vccd1 vccd1 _7623_/B sky130_fd_sc_hd__mux2_1
X_4834_ _4908_/A _4961_/A _5230_/A vssd1 vssd1 vccd1 vccd1 _4834_/X sky130_fd_sc_hd__o21a_1
X_7553_ _8721_/Q vssd1 vssd1 vccd1 vccd1 _8539_/A sky130_fd_sc_hd__clkbuf_2
X_4765_ _4803_/B _4765_/B vssd1 vssd1 vccd1 vccd1 _4766_/C sky130_fd_sc_hd__nand2_1
X_6504_ _6539_/A _6502_/X _6533_/A _8694_/Q vssd1 vssd1 vccd1 vccd1 _6505_/B sky130_fd_sc_hd__a31oi_1
X_7484_ _7480_/A _7480_/B _7480_/C _7367_/A vssd1 vssd1 vccd1 vccd1 _7485_/A sky130_fd_sc_hd__a31o_1
X_4696_ _5259_/A _4695_/A _4695_/Y _4677_/X vssd1 vssd1 vccd1 vccd1 _8595_/D sky130_fd_sc_hd__o211a_1
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6435_ _6435_/A _6435_/B vssd1 vssd1 vccd1 vccd1 _8673_/D sky130_fd_sc_hd__nor2_1
X_6366_ _6367_/A _6367_/B _6367_/C vssd1 vssd1 vccd1 vccd1 _6366_/Y sky130_fd_sc_hd__o21ai_1
X_8105_ _8042_/B _8105_/B vssd1 vssd1 vccd1 vccd1 _8105_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5317_ _6478_/A _5374_/A _5317_/C vssd1 vssd1 vccd1 vccd1 _5318_/A sky130_fd_sc_hd__and3_1
X_8036_ _8218_/A _7962_/B _7966_/B _7964_/X vssd1 vssd1 vccd1 vccd1 _8038_/B sky130_fd_sc_hd__a31oi_1
X_6297_ _6297_/A _6297_/B vssd1 vssd1 vccd1 vccd1 _6298_/B sky130_fd_sc_hd__xnor2_4
X_5248_ _5248_/A _5248_/B _5248_/C _5248_/D vssd1 vssd1 vccd1 vccd1 _5248_/X sky130_fd_sc_hd__or4_1
XFILLER_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5179_ _4728_/A _5170_/X _5178_/X _4701_/A vssd1 vssd1 vccd1 vccd1 _5179_/X sky130_fd_sc_hd__a211o_1
XFILLER_28_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8869_ _8869_/A _4386_/Y vssd1 vssd1 vccd1 vccd1 io_out[16] sky130_fd_sc_hd__ebufn_8
XFILLER_101_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4550_ _8615_/Q _4552_/B vssd1 vssd1 vccd1 vccd1 _4551_/A sky130_fd_sc_hd__and2_1
X_4481_ _4824_/B vssd1 vssd1 vccd1 vccd1 _4850_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6220_ _5996_/B _6220_/B vssd1 vssd1 vccd1 vccd1 _6220_/X sky130_fd_sc_hd__and2b_1
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6151_ _6151_/A _6151_/B vssd1 vssd1 vccd1 vccd1 _6151_/Y sky130_fd_sc_hd__nand2_1
XFILLER_97_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5102_ _5180_/A _5252_/A _5102_/C vssd1 vssd1 vccd1 vccd1 _5103_/B sky130_fd_sc_hd__or3_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6082_ _6214_/A _6082_/B vssd1 vssd1 vccd1 vccd1 _6083_/C sky130_fd_sc_hd__nand2_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5033_ _5190_/B _5024_/X _5020_/X _5028_/X _5032_/X vssd1 vssd1 vccd1 vccd1 _5034_/B
+ sky130_fd_sc_hd__o32a_1
XFILLER_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6984_ _6999_/A _6999_/B vssd1 vssd1 vccd1 vccd1 _6985_/B sky130_fd_sc_hd__xnor2_1
XFILLER_80_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8723_ input3/X _8723_/D vssd1 vssd1 vccd1 vccd1 _8723_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5935_ _5935_/A _5935_/B _5935_/C vssd1 vssd1 vccd1 vccd1 _5936_/B sky130_fd_sc_hd__nor3_1
XFILLER_25_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5866_ _5859_/A _5859_/B _5865_/X vssd1 vssd1 vccd1 vccd1 _5943_/A sky130_fd_sc_hd__a21oi_1
X_8654_ input3/X _8654_/D vssd1 vssd1 vccd1 vccd1 _8654_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7605_ _7604_/Y _7583_/X _4650_/A vssd1 vssd1 vccd1 vccd1 _7605_/Y sky130_fd_sc_hd__a21oi_1
X_4817_ _4865_/B vssd1 vssd1 vccd1 vccd1 _4859_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_33_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8585_ input3/X _8585_/D vssd1 vssd1 vccd1 vccd1 _8585_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5797_ _5726_/A _5809_/A _5727_/B _5731_/A vssd1 vssd1 vccd1 vccd1 _5812_/A sky130_fd_sc_hd__a22o_1
X_7536_ _7537_/A _7537_/B vssd1 vssd1 vccd1 vccd1 _7543_/B sky130_fd_sc_hd__nand2_1
X_4748_ _4745_/Y _4747_/X _4784_/A vssd1 vssd1 vccd1 vccd1 _8604_/D sky130_fd_sc_hd__a21oi_1
X_7467_ _7467_/A _7467_/B vssd1 vssd1 vccd1 vccd1 _7467_/X sky130_fd_sc_hd__or2_1
X_4679_ _5243_/A vssd1 vssd1 vccd1 vccd1 _4970_/A sky130_fd_sc_hd__buf_2
X_8729__7 vssd1 vssd1 vccd1 vccd1 _8729__7/HI _8824_/A sky130_fd_sc_hd__conb_1
X_6418_ _6418_/A vssd1 vssd1 vccd1 vccd1 _8668_/D sky130_fd_sc_hd__clkbuf_1
X_7398_ _7398_/A _7398_/B vssd1 vssd1 vccd1 vccd1 _7399_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6349_ _6346_/A _5412_/X _5413_/X _6348_/Y vssd1 vssd1 vccd1 vccd1 _8659_/D sky130_fd_sc_hd__a22o_1
XFILLER_88_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8019_ _8019_/A _8019_/B vssd1 vssd1 vccd1 vccd1 _8099_/B sky130_fd_sc_hd__nand2_1
XFILLER_48_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5720_ _5721_/A _5721_/B vssd1 vssd1 vccd1 vccd1 _5720_/X sky130_fd_sc_hd__or2_1
X_5651_ _6323_/C _6123_/A _5959_/A _5650_/Y vssd1 vssd1 vccd1 vccd1 _5697_/A sky130_fd_sc_hd__o31a_1
X_8370_ _8370_/A _8370_/B vssd1 vssd1 vccd1 vccd1 _8371_/B sky130_fd_sc_hd__xnor2_1
X_5582_ _5731_/A _5582_/B vssd1 vssd1 vccd1 vccd1 _5721_/B sky130_fd_sc_hd__xor2_1
X_4602_ _8576_/Q _4604_/C _4595_/X vssd1 vssd1 vccd1 vccd1 _4603_/B sky130_fd_sc_hd__o21ai_1
X_7321_ _7326_/A _7326_/B _7321_/C vssd1 vssd1 vccd1 vccd1 _7323_/B sky130_fd_sc_hd__nand3_1
X_4533_ _6777_/B _4533_/B vssd1 vssd1 vccd1 vccd1 _4662_/B sky130_fd_sc_hd__nor2_1
X_7252_ _7317_/A _7317_/B vssd1 vssd1 vccd1 vccd1 _7252_/Y sky130_fd_sc_hd__nand2_1
XFILLER_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6203_ _6203_/A _6203_/B vssd1 vssd1 vccd1 vccd1 _6204_/B sky130_fd_sc_hd__and2_1
X_4464_ _6556_/B vssd1 vssd1 vccd1 vccd1 _4662_/A sky130_fd_sc_hd__clkbuf_2
X_4395_ _4395_/A vssd1 vssd1 vccd1 vccd1 _4395_/Y sky130_fd_sc_hd__inv_2
X_7183_ _7254_/A _7254_/B _7182_/Y vssd1 vssd1 vccd1 vccd1 _7187_/A sky130_fd_sc_hd__a21o_1
X_6134_ _6134_/A _6134_/B vssd1 vssd1 vccd1 vccd1 _6135_/C sky130_fd_sc_hd__and2_1
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6065_ _6065_/A _6069_/B vssd1 vssd1 vccd1 vccd1 _6097_/B sky130_fd_sc_hd__xnor2_2
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5016_ _5245_/B _5231_/B _5102_/C _5057_/C vssd1 vssd1 vccd1 vccd1 _5168_/A sky130_fd_sc_hd__or4_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6967_ _6964_/Y _6965_/X _6824_/A _6895_/X vssd1 vssd1 vccd1 vccd1 _6988_/B sky130_fd_sc_hd__o211a_1
X_8706_ input3/X _8706_/D vssd1 vssd1 vccd1 vccd1 _8706_/Q sky130_fd_sc_hd__dfxtp_1
X_5918_ _5918_/A _5918_/B vssd1 vssd1 vccd1 vccd1 _5946_/B sky130_fd_sc_hd__xnor2_1
X_6898_ _7023_/A vssd1 vssd1 vccd1 vccd1 _7131_/A sky130_fd_sc_hd__clkbuf_2
X_5849_ _6203_/A _5849_/B vssd1 vssd1 vccd1 vccd1 _5850_/C sky130_fd_sc_hd__nor2_1
XFILLER_42_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8637_ input3/X _8637_/D vssd1 vssd1 vccd1 vccd1 _8637_/Q sky130_fd_sc_hd__dfxtp_1
X_8568_ _8568_/A _8568_/B vssd1 vssd1 vccd1 vccd1 _8568_/Y sky130_fd_sc_hd__nor2_1
X_7519_ _7518_/B _7525_/A vssd1 vssd1 vccd1 vccd1 _7520_/B sky130_fd_sc_hd__and2b_1
X_8499_ _8499_/A _8499_/B vssd1 vssd1 vccd1 vccd1 _8502_/A sky130_fd_sc_hd__xor2_1
XFILLER_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7870_ _8317_/A _8326_/A vssd1 vssd1 vccd1 vccd1 _7879_/A sky130_fd_sc_hd__nor2_1
X_6821_ _6897_/A _6897_/B vssd1 vssd1 vccd1 vccd1 _6823_/C sky130_fd_sc_hd__xnor2_1
XFILLER_23_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6752_ _6768_/B _6769_/C vssd1 vssd1 vccd1 vccd1 _7184_/A sky130_fd_sc_hd__xor2_2
X_6683_ _6799_/A vssd1 vssd1 vccd1 vccd1 _6919_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5703_ _5704_/A _5704_/B vssd1 vssd1 vccd1 vccd1 _6063_/B sky130_fd_sc_hd__nor2_1
X_8422_ _8482_/A _8482_/B vssd1 vssd1 vccd1 vccd1 _8423_/B sky130_fd_sc_hd__xnor2_1
X_5634_ _5647_/A _5647_/B vssd1 vssd1 vccd1 vccd1 _5666_/A sky130_fd_sc_hd__xnor2_2
X_8353_ _8297_/A _8353_/B vssd1 vssd1 vccd1 vccd1 _8353_/X sky130_fd_sc_hd__and2b_1
X_7304_ _7327_/A _7327_/B _7303_/Y vssd1 vssd1 vccd1 vccd1 _7310_/A sky130_fd_sc_hd__o21a_1
X_5565_ _5600_/A _5565_/B vssd1 vssd1 vccd1 vccd1 _5567_/C sky130_fd_sc_hd__and2_1
X_8284_ _8054_/A _8360_/A _8284_/C vssd1 vssd1 vccd1 vccd1 _8360_/B sky130_fd_sc_hd__nand3b_1
X_4516_ _4516_/A vssd1 vssd1 vccd1 vccd1 _8865_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5496_ _8658_/Q vssd1 vssd1 vccd1 vccd1 _6343_/S sky130_fd_sc_hd__inv_2
X_4447_ _4450_/A vssd1 vssd1 vccd1 vccd1 _4447_/Y sky130_fd_sc_hd__inv_2
X_7235_ _7308_/A _7234_/X _7200_/Y vssd1 vssd1 vccd1 vccd1 _7341_/B sky130_fd_sc_hd__o21a_1
X_7166_ _7293_/A _7246_/B vssd1 vssd1 vccd1 vccd1 _7168_/A sky130_fd_sc_hd__nand2_1
XFILLER_98_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4378_ _4396_/A vssd1 vssd1 vccd1 vccd1 _4383_/A sky130_fd_sc_hd__buf_6
X_6117_ _6117_/A _6117_/B vssd1 vssd1 vccd1 vccd1 _6121_/A sky130_fd_sc_hd__or2_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7097_ _7068_/A _7068_/B _7072_/A vssd1 vssd1 vccd1 vccd1 _7100_/A sky130_fd_sc_hd__a21bo_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6048_ _6054_/A _6054_/B vssd1 vssd1 vccd1 vccd1 _6077_/A sky130_fd_sc_hd__xor2_1
XFILLER_81_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7999_ _7923_/A _7923_/B _7998_/Y vssd1 vssd1 vccd1 vccd1 _8000_/B sky130_fd_sc_hd__o21ai_1
XFILLER_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8808__86 vssd1 vssd1 vccd1 vccd1 _8808__86/HI _8917_/A sky130_fd_sc_hd__conb_1
XFILLER_76_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5350_ _6471_/C _5352_/C _5374_/A vssd1 vssd1 vccd1 vccd1 _5350_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_99_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5281_ _8657_/Q _5271_/X _5280_/X _5273_/X vssd1 vssd1 vccd1 vccd1 _8615_/D sky130_fd_sc_hd__o211a_1
X_7020_ _7020_/A _7065_/B vssd1 vssd1 vccd1 vccd1 _7133_/A sky130_fd_sc_hd__or2b_1
XFILLER_4_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7922_ _7985_/C _7922_/B vssd1 vssd1 vccd1 vccd1 _7923_/B sky130_fd_sc_hd__xnor2_1
XFILLER_55_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7853_ _8205_/A _7853_/B _7853_/C vssd1 vssd1 vccd1 vccd1 _7853_/X sky130_fd_sc_hd__and3_1
XFILLER_23_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6804_ _6804_/A _6804_/B vssd1 vssd1 vccd1 vccd1 _6897_/A sky130_fd_sc_hd__xor2_2
X_7784_ _8060_/A _7784_/B vssd1 vssd1 vccd1 vccd1 _7786_/A sky130_fd_sc_hd__and2_1
X_4996_ _5023_/A _5086_/A _5167_/B vssd1 vssd1 vccd1 vccd1 _5135_/D sky130_fd_sc_hd__nor3_1
X_6735_ _6735_/A _6735_/B vssd1 vssd1 vccd1 vccd1 _7190_/A sky130_fd_sc_hd__nor2_1
XFILLER_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6666_ _6660_/A _6652_/B _6624_/B _6665_/X vssd1 vssd1 vccd1 vccd1 _6674_/B sky130_fd_sc_hd__a31o_1
X_8405_ _8327_/A _8407_/S _8328_/B _8331_/B vssd1 vssd1 vccd1 vccd1 _8408_/A sky130_fd_sc_hd__a22o_1
X_6597_ _7505_/A vssd1 vssd1 vccd1 vccd1 _7493_/A sky130_fd_sc_hd__inv_2
X_5617_ _5617_/A _8652_/Q vssd1 vssd1 vccd1 vccd1 _5617_/X sky130_fd_sc_hd__or2b_1
X_8336_ _8410_/A _8337_/B _8409_/B vssd1 vssd1 vccd1 vccd1 _8415_/A sky130_fd_sc_hd__a21o_1
X_5548_ _6009_/A _5561_/A vssd1 vssd1 vccd1 vccd1 _5898_/A sky130_fd_sc_hd__or2_2
X_8267_ _8267_/A _8267_/B vssd1 vssd1 vccd1 vccd1 _8497_/B sky130_fd_sc_hd__nor2_1
X_7218_ _7462_/A _7218_/B vssd1 vssd1 vccd1 vccd1 _7287_/A sky130_fd_sc_hd__xnor2_1
X_5479_ _5539_/B vssd1 vssd1 vccd1 vccd1 _5801_/C sky130_fd_sc_hd__buf_2
X_8198_ _8385_/A _8199_/B vssd1 vssd1 vccd1 vccd1 _8313_/A sky130_fd_sc_hd__nor2_1
XFILLER_48_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7149_ _7015_/B _7149_/B vssd1 vssd1 vccd1 vccd1 _7149_/X sky130_fd_sc_hd__and2b_1
XFILLER_58_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4850_ _4850_/A _4850_/B _5026_/A _4849_/A vssd1 vssd1 vccd1 vccd1 _5010_/B sky130_fd_sc_hd__or4b_2
XFILLER_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4781_ _4781_/A _4781_/B _5227_/A vssd1 vssd1 vccd1 vccd1 _4782_/B sky130_fd_sc_hd__and3_1
X_6520_ _6520_/A _6526_/B vssd1 vssd1 vccd1 vccd1 _6521_/B sky130_fd_sc_hd__and2_1
XFILLER_9_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6451_ _6450_/B _8677_/Q _6445_/B _8679_/Q vssd1 vssd1 vccd1 vccd1 _6452_/C sky130_fd_sc_hd__a31o_1
X_5402_ _5441_/A _5447_/A _5402_/C _5402_/D vssd1 vssd1 vccd1 vccd1 _5403_/B sky130_fd_sc_hd__or4_1
X_6382_ _8675_/Q vssd1 vssd1 vccd1 vccd1 _6441_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_8121_ _8214_/A _8214_/B vssd1 vssd1 vccd1 vccd1 _8132_/A sky130_fd_sc_hd__xnor2_2
X_5333_ _5333_/A vssd1 vssd1 vccd1 vccd1 _8629_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8052_ _8196_/A _8363_/A vssd1 vssd1 vccd1 vccd1 _8054_/B sky130_fd_sc_hd__xnor2_1
X_5264_ _5259_/B _4681_/B _4709_/A _5259_/A vssd1 vssd1 vccd1 vccd1 _5265_/C sky130_fd_sc_hd__o211a_1
X_7003_ _6980_/A _6979_/B _6979_/A vssd1 vssd1 vccd1 vccd1 _7012_/A sky130_fd_sc_hd__a21oi_2
X_5195_ _5245_/A _5199_/A _5194_/X vssd1 vssd1 vccd1 vccd1 _5195_/Y sky130_fd_sc_hd__a21oi_1
X_8799__77 vssd1 vssd1 vccd1 vccd1 _8799__77/HI _8908_/A sky130_fd_sc_hd__conb_1
XFILLER_95_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8885_ _8885_/A _4406_/Y vssd1 vssd1 vccd1 vccd1 io_out[32] sky130_fd_sc_hd__ebufn_8
X_7905_ _7796_/B _7792_/B _7904_/X vssd1 vssd1 vccd1 vccd1 _7916_/A sky130_fd_sc_hd__a21oi_1
XFILLER_24_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7836_ _7904_/A _7836_/B _7836_/C vssd1 vssd1 vccd1 vccd1 _8508_/A sky130_fd_sc_hd__and3_1
XFILLER_34_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7767_ _7766_/A _7766_/C _7766_/B vssd1 vssd1 vccd1 vccd1 _7957_/D sky130_fd_sc_hd__a21oi_2
XFILLER_11_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4979_ _4979_/A _5145_/B vssd1 vssd1 vccd1 vccd1 _5055_/B sky130_fd_sc_hd__or2_1
X_7698_ _7722_/A _7722_/B _7697_/X vssd1 vssd1 vccd1 vccd1 _7745_/B sky130_fd_sc_hd__a21o_2
X_6718_ _7293_/B _6717_/X _6718_/S vssd1 vssd1 vccd1 vccd1 _6814_/A sky130_fd_sc_hd__mux2_4
X_6649_ _6831_/B _6709_/B vssd1 vssd1 vccd1 vccd1 _6651_/B sky130_fd_sc_hd__xnor2_2
X_8319_ _8319_/A _8319_/B _8319_/C vssd1 vssd1 vccd1 vccd1 _8320_/B sky130_fd_sc_hd__nor3_1
XFILLER_3_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5951_ _6277_/A _5951_/B vssd1 vssd1 vccd1 vccd1 _5951_/Y sky130_fd_sc_hd__nor2_1
XFILLER_18_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4902_ _5193_/A vssd1 vssd1 vccd1 vccd1 _5098_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_8670_ input3/X _8670_/D vssd1 vssd1 vccd1 vccd1 _8670_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5882_ _5882_/A _5882_/B vssd1 vssd1 vccd1 vccd1 _6143_/B sky130_fd_sc_hd__nor2_1
X_7621_ _8712_/Q _7621_/B vssd1 vssd1 vccd1 vccd1 _7621_/X sky130_fd_sc_hd__or2_1
X_4833_ _5119_/A _5248_/A _4832_/X vssd1 vssd1 vccd1 vccd1 _5230_/A sky130_fd_sc_hd__nor3b_1
XFILLER_21_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7552_ _7552_/A vssd1 vssd1 vccd1 vccd1 _7552_/Y sky130_fd_sc_hd__inv_2
X_4764_ _4803_/B _4765_/B vssd1 vssd1 vccd1 vccd1 _4775_/C sky130_fd_sc_hd__nor2_1
X_7483_ _7480_/X _7481_/Y _7482_/Y _7477_/B vssd1 vssd1 vccd1 vccd1 _7486_/B sky130_fd_sc_hd__a2bb2o_1
X_6503_ _6536_/A _6531_/B vssd1 vssd1 vccd1 vccd1 _6533_/A sky130_fd_sc_hd__or2_1
X_4695_ _4695_/A _5251_/A vssd1 vssd1 vccd1 vccd1 _4695_/Y sky130_fd_sc_hd__nand2_1
X_6434_ _8673_/Q _6436_/C _6427_/X vssd1 vssd1 vccd1 vccd1 _6435_/B sky130_fd_sc_hd__o21ai_1
X_6365_ _6358_/B _6359_/Y _5384_/Y vssd1 vssd1 vccd1 vccd1 _6367_/C sky130_fd_sc_hd__o21ai_1
X_8104_ _8072_/A _8072_/B _8103_/Y vssd1 vssd1 vccd1 vccd1 _8189_/A sky130_fd_sc_hd__a21boi_1
X_6296_ _6296_/A _6296_/B vssd1 vssd1 vccd1 vccd1 _6297_/B sky130_fd_sc_hd__xnor2_2
X_5316_ _8625_/Q _8624_/Q vssd1 vssd1 vccd1 vccd1 _5317_/C sky130_fd_sc_hd__nand2_1
XFILLER_88_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8035_ _7972_/A _8317_/B _7973_/B _8321_/A vssd1 vssd1 vccd1 vccd1 _8040_/A sky130_fd_sc_hd__a2bb2o_1
X_5247_ _5256_/B _5115_/X _5054_/D _5103_/X _4969_/B vssd1 vssd1 vccd1 vccd1 _5248_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_29_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5178_ _5134_/X _5171_/X _5177_/X _4686_/A vssd1 vssd1 vccd1 vccd1 _5178_/X sky130_fd_sc_hd__o211a_1
XFILLER_29_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8868_ _8868_/A _4385_/Y vssd1 vssd1 vccd1 vccd1 io_out[15] sky130_fd_sc_hd__ebufn_8
XFILLER_101_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7819_ _7819_/A _7819_/B vssd1 vssd1 vccd1 vccd1 _7820_/B sky130_fd_sc_hd__and2_1
XFILLER_12_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4480_ _4831_/B vssd1 vssd1 vccd1 vccd1 _4824_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6150_ _6096_/A _6095_/B _6095_/C vssd1 vssd1 vccd1 vccd1 _6151_/B sky130_fd_sc_hd__o21ai_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5101_ _5101_/A vssd1 vssd1 vccd1 vccd1 _5252_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6081_ _6081_/A _6081_/B vssd1 vssd1 vccd1 vccd1 _6085_/A sky130_fd_sc_hd__xnor2_1
XFILLER_97_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5032_ _5190_/B _5029_/X _5030_/X _5072_/C vssd1 vssd1 vccd1 vccd1 _5032_/X sky130_fd_sc_hd__o22a_1
X_8769__47 vssd1 vssd1 vccd1 vccd1 _8769__47/HI _8878_/A sky130_fd_sc_hd__conb_1
XFILLER_65_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6983_ _6887_/A _6886_/B _6886_/A vssd1 vssd1 vccd1 vccd1 _6999_/B sky130_fd_sc_hd__a21boi_1
XFILLER_65_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8722_ input3/X _8722_/D vssd1 vssd1 vccd1 vccd1 _8722_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5934_ _5935_/A _5935_/B _5935_/C vssd1 vssd1 vccd1 vccd1 _5936_/A sky130_fd_sc_hd__o21a_1
X_5865_ _5845_/A _5865_/B vssd1 vssd1 vccd1 vccd1 _5865_/X sky130_fd_sc_hd__and2b_1
X_8653_ input3/X _8653_/D vssd1 vssd1 vccd1 vccd1 _8653_/Q sky130_fd_sc_hd__dfxtp_1
X_7604_ _7604_/A vssd1 vssd1 vccd1 vccd1 _7604_/Y sky130_fd_sc_hd__inv_2
X_4816_ _4839_/A vssd1 vssd1 vccd1 vccd1 _4865_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_8584_ input3/X _8584_/D vssd1 vssd1 vccd1 vccd1 _8584_/Q sky130_fd_sc_hd__dfxtp_1
X_5796_ _6005_/A _5896_/B vssd1 vssd1 vccd1 vccd1 _5805_/A sky130_fd_sc_hd__xnor2_1
X_4747_ _4745_/A _4822_/A _4746_/Y vssd1 vssd1 vccd1 vccd1 _4747_/X sky130_fd_sc_hd__a21o_1
XFILLER_31_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7535_ _7533_/A _7537_/B _7543_/A vssd1 vssd1 vccd1 vccd1 _7539_/A sky130_fd_sc_hd__o21ai_1
X_7466_ _7467_/A _7467_/B _7488_/A vssd1 vssd1 vccd1 vccd1 _7466_/X sky130_fd_sc_hd__a21o_1
X_4678_ _4661_/A _4739_/A _4697_/B _4677_/X vssd1 vssd1 vccd1 vccd1 _8592_/D sky130_fd_sc_hd__o211a_1
X_7397_ _7397_/A _7397_/B vssd1 vssd1 vccd1 vccd1 _7416_/B sky130_fd_sc_hd__xnor2_1
X_6417_ _6422_/C _6417_/B _6461_/B vssd1 vssd1 vccd1 vccd1 _6418_/A sky130_fd_sc_hd__and3b_1
X_6348_ _8658_/Q _6348_/B vssd1 vssd1 vccd1 vccd1 _6348_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6279_ _6188_/A _6279_/B vssd1 vssd1 vccd1 vccd1 _6279_/X sky130_fd_sc_hd__and2b_1
XFILLER_102_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8018_ _8018_/A _8018_/B vssd1 vssd1 vccd1 vccd1 _8090_/A sky130_fd_sc_hd__and2_1
XFILLER_91_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8783__61 vssd1 vssd1 vccd1 vccd1 _8783__61/HI _8892_/A sky130_fd_sc_hd__conb_1
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5650_ _5701_/A _5695_/B vssd1 vssd1 vccd1 vccd1 _5650_/Y sky130_fd_sc_hd__nand2_1
XFILLER_43_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4601_ _8576_/Q _4604_/C vssd1 vssd1 vccd1 vccd1 _4603_/A sky130_fd_sc_hd__and2_1
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5581_ _5801_/C _5906_/A _5589_/A _5595_/A vssd1 vssd1 vccd1 vccd1 _5582_/B sky130_fd_sc_hd__o22a_1
X_7320_ _7320_/A _7320_/B vssd1 vssd1 vccd1 vccd1 _7321_/C sky130_fd_sc_hd__xor2_1
XFILLER_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4532_ _8599_/Q vssd1 vssd1 vccd1 vccd1 _6777_/B sky130_fd_sc_hd__clkbuf_2
X_7251_ _7315_/A _7251_/B vssd1 vssd1 vccd1 vccd1 _7318_/B sky130_fd_sc_hd__xor2_2
X_4463_ _8596_/Q vssd1 vssd1 vccd1 vccd1 _6556_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_89_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6202_ _6202_/A _5998_/A vssd1 vssd1 vccd1 vccd1 _6207_/A sky130_fd_sc_hd__or2b_1
X_4394_ _4395_/A vssd1 vssd1 vccd1 vccd1 _4394_/Y sky130_fd_sc_hd__inv_2
X_7182_ _7182_/A _7182_/B vssd1 vssd1 vccd1 vccd1 _7182_/Y sky130_fd_sc_hd__nor2_1
X_6133_ _6046_/Y _6108_/A _6117_/A vssd1 vssd1 vccd1 vccd1 _6138_/A sky130_fd_sc_hd__o21ba_1
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6064_ _5781_/A _6063_/Y _5706_/A _5706_/B vssd1 vssd1 vccd1 vccd1 _6069_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5015_ _5015_/A vssd1 vssd1 vccd1 vccd1 _5245_/B sky130_fd_sc_hd__clkbuf_2
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6966_ _6824_/A _6895_/X _6964_/Y _6965_/X vssd1 vssd1 vccd1 vccd1 _6998_/A sky130_fd_sc_hd__a211oi_2
XFILLER_53_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5917_ _5917_/A _5977_/B vssd1 vssd1 vccd1 vccd1 _5918_/B sky130_fd_sc_hd__xnor2_1
X_8705_ input3/X _8705_/D vssd1 vssd1 vccd1 vccd1 _8705_/Q sky130_fd_sc_hd__dfxtp_1
X_8731__9 vssd1 vssd1 vccd1 vccd1 _8731__9/HI _8826_/A sky130_fd_sc_hd__conb_1
X_6897_ _6897_/A _6897_/B vssd1 vssd1 vccd1 vccd1 _6897_/Y sky130_fd_sc_hd__nand2_1
XFILLER_42_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8636_ input3/X _8636_/D vssd1 vssd1 vccd1 vccd1 _8636_/Q sky130_fd_sc_hd__dfxtp_1
X_5848_ _5956_/A vssd1 vssd1 vccd1 vccd1 _6203_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_8567_ _8566_/X _8562_/A _8567_/S vssd1 vssd1 vccd1 vccd1 _8568_/B sky130_fd_sc_hd__mux2_1
X_5779_ _5937_/A _5779_/B vssd1 vssd1 vccd1 vccd1 _5781_/B sky130_fd_sc_hd__nor2_1
X_7518_ _7525_/A _7518_/B vssd1 vssd1 vccd1 vccd1 _7520_/A sky130_fd_sc_hd__and2b_1
X_8498_ _8497_/B _8497_/C _8497_/A vssd1 vssd1 vccd1 vccd1 _8498_/X sky130_fd_sc_hd__o21a_1
X_7449_ _7449_/A _7449_/B _7449_/C vssd1 vssd1 vccd1 vccd1 _7449_/X sky130_fd_sc_hd__and3_1
XFILLER_89_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8739__17 vssd1 vssd1 vccd1 vccd1 _8739__17/HI _8834_/A sky130_fd_sc_hd__conb_1
XFILLER_75_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6820_ _6896_/A _6820_/B vssd1 vssd1 vccd1 vccd1 _6897_/B sky130_fd_sc_hd__xnor2_1
XFILLER_35_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6751_ _6751_/A _7179_/A vssd1 vssd1 vccd1 vccd1 _6769_/C sky130_fd_sc_hd__xnor2_2
X_6682_ _6656_/B _6657_/B _6657_/C _6629_/A vssd1 vssd1 vccd1 vccd1 _6799_/A sky130_fd_sc_hd__a31o_1
X_5702_ _6044_/A _5956_/A _6049_/B _6107_/B _6180_/A vssd1 vssd1 vccd1 vccd1 _5704_/B
+ sky130_fd_sc_hd__o32a_1
X_8421_ _8421_/A _8421_/B vssd1 vssd1 vccd1 vccd1 _8482_/B sky130_fd_sc_hd__xor2_1
X_5633_ _5633_/A _5633_/B vssd1 vssd1 vccd1 vccd1 _5647_/B sky130_fd_sc_hd__nor2_2
XFILLER_31_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8352_ _8349_/A _8352_/B vssd1 vssd1 vccd1 vccd1 _8425_/B sky130_fd_sc_hd__and2b_1
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5564_ _6034_/A _5794_/B _5794_/C _6003_/A vssd1 vssd1 vccd1 vccd1 _5565_/B sky130_fd_sc_hd__a31o_1
X_7303_ _7398_/A _7303_/B vssd1 vssd1 vccd1 vccd1 _7303_/Y sky130_fd_sc_hd__nand2_1
X_4515_ _4745_/A _4781_/B _4542_/A _4541_/C vssd1 vssd1 vccd1 vccd1 _4516_/A sky130_fd_sc_hd__or4_2
X_8283_ _8283_/A _8305_/B vssd1 vssd1 vccd1 vccd1 _8360_/A sky130_fd_sc_hd__or2_1
X_5495_ _5794_/A _5558_/A vssd1 vssd1 vccd1 vccd1 _5511_/A sky130_fd_sc_hd__nand2_1
X_4446_ _4450_/A vssd1 vssd1 vccd1 vccd1 _4446_/Y sky130_fd_sc_hd__inv_2
X_7234_ _7234_/A _7234_/B vssd1 vssd1 vccd1 vccd1 _7234_/X sky130_fd_sc_hd__or2_1
X_4377_ _4377_/A vssd1 vssd1 vccd1 vccd1 _4377_/Y sky130_fd_sc_hd__inv_2
X_7165_ _7165_/A vssd1 vssd1 vccd1 vccd1 _7293_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_98_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6116_ _5954_/A _5701_/A _5953_/Y _6112_/X _6114_/X vssd1 vssd1 vccd1 vccd1 _6117_/B
+ sky130_fd_sc_hd__a2111oi_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7096_ _7096_/A _7096_/B vssd1 vssd1 vccd1 vccd1 _7113_/A sky130_fd_sc_hd__xnor2_1
XFILLER_58_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6047_ _5953_/B _6108_/A _6109_/B _6046_/Y vssd1 vssd1 vccd1 vccd1 _6054_/B sky130_fd_sc_hd__a211o_1
XFILLER_39_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7998_ _7998_/A _7998_/B vssd1 vssd1 vccd1 vccd1 _7998_/Y sky130_fd_sc_hd__nand2_1
X_8753__31 vssd1 vssd1 vccd1 vccd1 _8753__31/HI _8848_/A sky130_fd_sc_hd__conb_1
X_6949_ _6949_/A _7025_/B vssd1 vssd1 vccd1 vccd1 _6950_/B sky130_fd_sc_hd__xor2_2
XFILLER_22_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8619_ input3/X _8619_/D vssd1 vssd1 vccd1 vccd1 _8619_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5280_ _8615_/Q _5288_/B vssd1 vssd1 vccd1 vccd1 _5280_/X sky130_fd_sc_hd__or2_1
XFILLER_4_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7921_ _8006_/B _7921_/B vssd1 vssd1 vccd1 vccd1 _7922_/B sky130_fd_sc_hd__nor2_1
XFILLER_36_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7852_ _7775_/A _7852_/B vssd1 vssd1 vccd1 vccd1 _7948_/A sky130_fd_sc_hd__and2b_1
XFILLER_36_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6803_ _6803_/A _6803_/B vssd1 vssd1 vccd1 vccd1 _6804_/B sky130_fd_sc_hd__xor2_1
XFILLER_63_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7783_ _7783_/A _7574_/X vssd1 vssd1 vccd1 vccd1 _7784_/B sky130_fd_sc_hd__or2b_1
X_4995_ _4995_/A vssd1 vssd1 vccd1 vccd1 _5190_/A sky130_fd_sc_hd__clkbuf_2
X_6734_ _6734_/A _6734_/B _6734_/C vssd1 vssd1 vccd1 vccd1 _6735_/B sky130_fd_sc_hd__and3_1
XFILLER_23_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8404_ _8404_/A _8404_/B vssd1 vssd1 vccd1 vccd1 _8415_/B sky130_fd_sc_hd__nand2_1
X_6665_ _8692_/Q _7658_/B vssd1 vssd1 vccd1 vccd1 _6665_/X sky130_fd_sc_hd__and2b_1
X_6596_ _6596_/A _6596_/B vssd1 vssd1 vccd1 vccd1 _7505_/A sky130_fd_sc_hd__xnor2_2
X_5616_ _5759_/A _5616_/B vssd1 vssd1 vccd1 vccd1 _5660_/A sky130_fd_sc_hd__nand2_1
X_8335_ _8410_/B _8410_/C vssd1 vssd1 vccd1 vccd1 _8409_/B sky130_fd_sc_hd__xnor2_1
X_5547_ _5482_/A _5546_/X _5508_/X _5506_/A vssd1 vssd1 vccd1 vccd1 _5561_/A sky130_fd_sc_hd__a31o_1
X_8266_ _8503_/B _8503_/C _8495_/A _8503_/A vssd1 vssd1 vccd1 vccd1 _8492_/B sky130_fd_sc_hd__a211o_1
X_5478_ _5494_/A _5533_/B vssd1 vssd1 vccd1 vccd1 _5539_/B sky130_fd_sc_hd__or2_1
X_7217_ _7217_/A _7217_/B vssd1 vssd1 vccd1 vccd1 _7218_/B sky130_fd_sc_hd__nor2_1
X_4429_ _4432_/A vssd1 vssd1 vccd1 vccd1 _4429_/Y sky130_fd_sc_hd__inv_2
X_8197_ _8382_/A _8196_/X _8144_/Y vssd1 vssd1 vccd1 vccd1 _8199_/B sky130_fd_sc_hd__a21o_1
XFILLER_59_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7148_ _7086_/A _7086_/B _7147_/Y vssd1 vssd1 vccd1 vccd1 _7156_/A sky130_fd_sc_hd__o21a_1
XFILLER_48_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7079_ _7078_/B _7078_/C _7078_/A vssd1 vssd1 vccd1 vccd1 _7081_/B sky130_fd_sc_hd__o21a_1
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4780_ _4824_/C _4897_/A vssd1 vssd1 vccd1 vccd1 _5227_/A sky130_fd_sc_hd__nor2_1
XFILLER_33_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6450_ _8679_/Q _6450_/B _6450_/C vssd1 vssd1 vccd1 vccd1 _6454_/B sky130_fd_sc_hd__and3_1
X_5401_ _5421_/A _5414_/A _5428_/A vssd1 vssd1 vccd1 vccd1 _5402_/D sky130_fd_sc_hd__o21a_1
X_6381_ _8680_/Q _8682_/Q _8681_/Q _8679_/Q vssd1 vssd1 vccd1 vccd1 _6398_/A sky130_fd_sc_hd__and4bb_1
X_8120_ _8120_/A _8120_/B vssd1 vssd1 vccd1 vccd1 _8214_/B sky130_fd_sc_hd__xnor2_2
X_5332_ _5337_/C _5332_/B _5354_/B vssd1 vssd1 vccd1 vccd1 _5333_/A sky130_fd_sc_hd__and3b_1
X_8051_ _8051_/A _8152_/A vssd1 vssd1 vccd1 vccd1 _8363_/A sky130_fd_sc_hd__nand2_4
X_5263_ _5263_/A _5263_/B _4820_/B vssd1 vssd1 vccd1 vccd1 _5269_/B sky130_fd_sc_hd__or3b_1
X_7002_ _6963_/A _6963_/B _7001_/X vssd1 vssd1 vccd1 vccd1 _7142_/B sky130_fd_sc_hd__a21bo_1
X_5194_ _5194_/A _5241_/A _5193_/Y vssd1 vssd1 vccd1 vccd1 _5194_/X sky130_fd_sc_hd__or3b_1
XFILLER_95_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8884_ _8884_/A _4405_/Y vssd1 vssd1 vccd1 vccd1 io_out[31] sky130_fd_sc_hd__ebufn_8
X_7904_ _7904_/A _8056_/B _7904_/C vssd1 vssd1 vccd1 vccd1 _7904_/X sky130_fd_sc_hd__and3_1
X_7835_ _7986_/A _7988_/A vssd1 vssd1 vccd1 vccd1 _7836_/C sky130_fd_sc_hd__or2_1
XFILLER_51_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7766_ _7766_/A _7766_/B _7766_/C vssd1 vssd1 vccd1 vccd1 _7957_/C sky130_fd_sc_hd__and3_1
XFILLER_51_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4978_ _4988_/A vssd1 vssd1 vccd1 vccd1 _5132_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7697_ _8720_/Q _8596_/Q vssd1 vssd1 vccd1 vccd1 _7697_/X sky130_fd_sc_hd__and2b_1
X_6717_ _6614_/X _6642_/X _6643_/X _6671_/B _6798_/A vssd1 vssd1 vccd1 vccd1 _6717_/X
+ sky130_fd_sc_hd__a311o_1
X_6648_ _6641_/X _7065_/A _6730_/A vssd1 vssd1 vccd1 vccd1 _6709_/B sky130_fd_sc_hd__a21oi_2
X_8318_ _8319_/B _8319_/C _8319_/A vssd1 vssd1 vccd1 vccd1 _8320_/A sky130_fd_sc_hd__o21a_1
X_6579_ _7297_/A _6647_/A vssd1 vssd1 vccd1 vccd1 _7439_/A sky130_fd_sc_hd__or2_2
XFILLER_3_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8249_ _8079_/B _8174_/B _8172_/Y vssd1 vssd1 vccd1 vccd1 _8251_/B sky130_fd_sc_hd__a21o_1
XFILLER_78_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5950_ _5950_/A _5929_/B vssd1 vssd1 vccd1 vccd1 _5972_/B sky130_fd_sc_hd__or2b_1
XFILLER_92_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4901_ _5115_/B _5151_/B _5118_/C vssd1 vssd1 vccd1 vccd1 _4901_/X sky130_fd_sc_hd__or3_1
XFILLER_45_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7620_ _7616_/A _7581_/X _7619_/Y _7541_/X vssd1 vssd1 vccd1 vccd1 _8713_/D sky130_fd_sc_hd__a211o_1
X_5881_ _5881_/A _5881_/B vssd1 vssd1 vccd1 vccd1 _5882_/B sky130_fd_sc_hd__and2_1
XFILLER_60_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4832_ _4897_/A _4897_/B _4836_/B _4960_/A _4908_/A vssd1 vssd1 vccd1 vccd1 _4832_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_21_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7551_ _8725_/Q vssd1 vssd1 vccd1 vccd1 _7875_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_21_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4763_ _5620_/A vssd1 vssd1 vccd1 vccd1 _4803_/B sky130_fd_sc_hd__inv_2
X_7482_ _7482_/A _7482_/B vssd1 vssd1 vccd1 vccd1 _7482_/Y sky130_fd_sc_hd__nand2_1
X_4694_ _4694_/A vssd1 vssd1 vccd1 vccd1 _5251_/A sky130_fd_sc_hd__clkbuf_2
X_6502_ _6514_/A _8688_/Q _6531_/B _6520_/A _6526_/A vssd1 vssd1 vccd1 vccd1 _6502_/X
+ sky130_fd_sc_hd__a2111o_1
X_6433_ _8673_/Q _6436_/C vssd1 vssd1 vccd1 vccd1 _6435_/A sky130_fd_sc_hd__and2_1
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6364_ _6375_/A _6364_/B vssd1 vssd1 vccd1 vccd1 _6367_/B sky130_fd_sc_hd__and2_1
X_8103_ _8103_/A _8103_/B vssd1 vssd1 vccd1 vccd1 _8103_/Y sky130_fd_sc_hd__nand2_1
X_6295_ _6295_/A _6295_/B vssd1 vssd1 vccd1 vccd1 _6296_/B sky130_fd_sc_hd__xnor2_1
X_5315_ _5320_/A vssd1 vssd1 vccd1 vccd1 _5374_/A sky130_fd_sc_hd__clkbuf_2
X_8034_ _8406_/A vssd1 vssd1 vccd1 vccd1 _8321_/A sky130_fd_sc_hd__clkbuf_2
X_5246_ _5105_/X _5245_/B _5118_/D _5245_/X vssd1 vssd1 vccd1 vccd1 _5246_/X sky130_fd_sc_hd__o31a_1
XFILLER_102_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5177_ _5105_/X _5173_/X _5176_/X _5139_/A vssd1 vssd1 vccd1 vccd1 _5177_/X sky130_fd_sc_hd__a211o_1
XFILLER_71_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8867_ _8867_/A _4383_/Y vssd1 vssd1 vccd1 vccd1 io_out[14] sky130_fd_sc_hd__ebufn_8
X_7818_ _7986_/A _8050_/A vssd1 vssd1 vccd1 vccd1 _8284_/C sky130_fd_sc_hd__or2_1
X_7749_ _8725_/Q _8601_/Q vssd1 vssd1 vccd1 vccd1 _7751_/A sky130_fd_sc_hd__and2b_1
XFILLER_86_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6080_ _6087_/A _6087_/B _6094_/B vssd1 vssd1 vccd1 vccd1 _6157_/A sky130_fd_sc_hd__or3b_2
X_5100_ _4686_/A _5090_/X _5099_/X _4694_/A vssd1 vssd1 vccd1 vccd1 _5100_/X sky130_fd_sc_hd__a211o_1
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5031_ _5091_/A _5046_/A vssd1 vssd1 vccd1 vccd1 _5072_/C sky130_fd_sc_hd__or2_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6982_ _6982_/A _6982_/B vssd1 vssd1 vccd1 vccd1 _6999_/A sky130_fd_sc_hd__xnor2_1
X_8721_ input3/X _8721_/D vssd1 vssd1 vccd1 vccd1 _8721_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5933_ _5976_/A _5933_/B vssd1 vssd1 vccd1 vccd1 _5935_/C sky130_fd_sc_hd__and2b_1
X_5864_ _5858_/A _5858_/B _5857_/A vssd1 vssd1 vccd1 vccd1 _5941_/A sky130_fd_sc_hd__o21ai_1
X_8652_ input3/X _8652_/D vssd1 vssd1 vccd1 vccd1 _8652_/Q sky130_fd_sc_hd__dfxtp_1
X_7603_ _7603_/A _7603_/B vssd1 vssd1 vccd1 vccd1 _7603_/Y sky130_fd_sc_hd__nor2_1
X_4815_ _4848_/A _4848_/B vssd1 vssd1 vccd1 vccd1 _4839_/A sky130_fd_sc_hd__or2_1
XFILLER_21_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8583_ input3/X _8583_/D vssd1 vssd1 vccd1 vccd1 _8583_/Q sky130_fd_sc_hd__dfxtp_1
X_5795_ _5795_/A _5895_/B vssd1 vssd1 vccd1 vccd1 _5896_/B sky130_fd_sc_hd__xnor2_1
X_7534_ _6513_/A _7543_/A _7532_/X _7533_/Y vssd1 vssd1 vccd1 vccd1 _8703_/D sky130_fd_sc_hd__a31o_1
X_4746_ _4745_/A _4822_/A _4675_/B vssd1 vssd1 vccd1 vccd1 _4746_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_31_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7465_ _7488_/B vssd1 vssd1 vccd1 vccd1 _7465_/Y sky130_fd_sc_hd__inv_2
X_4677_ _4717_/A vssd1 vssd1 vccd1 vccd1 _4677_/X sky130_fd_sc_hd__clkbuf_2
X_7396_ _7396_/A _7396_/B vssd1 vssd1 vccd1 vccd1 _7452_/A sky130_fd_sc_hd__xnor2_1
X_6416_ _8668_/Q _6416_/B vssd1 vssd1 vccd1 vccd1 _6417_/B sky130_fd_sc_hd__or2_1
X_6347_ _6347_/A _6347_/B vssd1 vssd1 vccd1 vccd1 _6348_/B sky130_fd_sc_hd__nand2_1
XFILLER_88_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6278_ _6278_/A _6278_/B vssd1 vssd1 vccd1 vccd1 _6296_/A sky130_fd_sc_hd__xnor2_1
X_8017_ _8017_/A _8015_/B vssd1 vssd1 vccd1 vccd1 _8263_/A sky130_fd_sc_hd__or2b_1
X_5229_ _5252_/A _5004_/C _5229_/C _5229_/D vssd1 vssd1 vccd1 vccd1 _5230_/C sky130_fd_sc_hd__and4bb_1
XFILLER_56_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8919_ _8919_/A _4444_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[28] sky130_fd_sc_hd__ebufn_8
XFILLER_71_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4600_ _4604_/C _4600_/B vssd1 vssd1 vccd1 vccd1 _8575_/D sky130_fd_sc_hd__nor2_1
X_5580_ _6009_/A _5580_/B vssd1 vssd1 vccd1 vccd1 _5589_/A sky130_fd_sc_hd__nor2_1
X_4531_ _5149_/A _4728_/B _5253_/A _4662_/A vssd1 vssd1 vccd1 vccd1 _4534_/C sky130_fd_sc_hd__o31a_1
X_7250_ _7317_/A _7317_/B vssd1 vssd1 vccd1 vccd1 _7250_/X sky130_fd_sc_hd__or2_1
XFILLER_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4462_ _7689_/B vssd1 vssd1 vccd1 vccd1 _7688_/B sky130_fd_sc_hd__buf_2
X_6201_ _6269_/A _6201_/B vssd1 vssd1 vccd1 vccd1 _6209_/A sky130_fd_sc_hd__nor2_1
X_4393_ _4395_/A vssd1 vssd1 vccd1 vccd1 _4393_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7181_ _7182_/A _7182_/B vssd1 vssd1 vccd1 vccd1 _7254_/B sky130_fd_sc_hd__xor2_1
X_6132_ _6142_/A _6142_/B vssd1 vssd1 vccd1 vccd1 _6140_/C sky130_fd_sc_hd__and2b_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6063_ _6063_/A _6063_/B vssd1 vssd1 vccd1 vccd1 _6063_/Y sky130_fd_sc_hd__nor2_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5014_ _5182_/C _5047_/B _5014_/C _5014_/D vssd1 vssd1 vccd1 vccd1 _5014_/X sky130_fd_sc_hd__or4_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6965_ _6964_/A _6964_/B _6964_/C vssd1 vssd1 vccd1 vccd1 _6965_/X sky130_fd_sc_hd__o21a_1
XFILLER_26_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8704_ input3/X _8704_/D vssd1 vssd1 vccd1 vccd1 _8704_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5916_ _5916_/A _5916_/B vssd1 vssd1 vccd1 vccd1 _5977_/B sky130_fd_sc_hd__xor2_1
XFILLER_41_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6896_ _6896_/A _6820_/B vssd1 vssd1 vccd1 vccd1 _6896_/X sky130_fd_sc_hd__or2b_1
X_8635_ input3/X _8635_/D vssd1 vssd1 vccd1 vccd1 _8635_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5847_ _6193_/A _5921_/B vssd1 vssd1 vccd1 vccd1 _5850_/B sky130_fd_sc_hd__xor2_1
XFILLER_21_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8566_ _8566_/A _8566_/B vssd1 vssd1 vccd1 vccd1 _8566_/X sky130_fd_sc_hd__or2_1
X_5778_ _5777_/A _5777_/B _5777_/C vssd1 vssd1 vccd1 vccd1 _5779_/B sky130_fd_sc_hd__a21oi_1
XFILLER_21_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8497_ _8497_/A _8497_/B _8497_/C vssd1 vssd1 vccd1 vccd1 _8497_/Y sky130_fd_sc_hd__nor3_1
X_4729_ _8593_/Q vssd1 vssd1 vccd1 vccd1 _5135_/A sky130_fd_sc_hd__clkbuf_2
X_7517_ _7514_/A _6511_/X _6513_/X _7516_/Y vssd1 vssd1 vccd1 vccd1 _8700_/D sky130_fd_sc_hd__a22o_1
X_7448_ _7436_/A _7436_/B _7446_/B _7447_/X vssd1 vssd1 vccd1 vccd1 _7474_/B sky130_fd_sc_hd__a31o_1
XFILLER_89_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7379_ _7385_/A _7385_/B vssd1 vssd1 vccd1 vccd1 _7380_/B sky130_fd_sc_hd__xor2_1
XFILLER_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6750_ _6947_/A vssd1 vssd1 vccd1 vccd1 _7179_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_63_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5701_ _5701_/A _5749_/B vssd1 vssd1 vccd1 vccd1 _6049_/B sky130_fd_sc_hd__xnor2_1
X_6681_ _6676_/X _6724_/A _6724_/B vssd1 vssd1 vccd1 vccd1 _6692_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8420_ _8435_/A _8435_/B vssd1 vssd1 vccd1 vccd1 _8421_/B sky130_fd_sc_hd__xor2_1
X_5632_ _5617_/A _8652_/Q vssd1 vssd1 vccd1 vccd1 _5633_/A sky130_fd_sc_hd__and2b_1
XFILLER_31_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8351_ _8348_/B _8351_/B vssd1 vssd1 vccd1 vccd1 _8425_/A sky130_fd_sc_hd__and2b_1
X_5563_ _5563_/A _5595_/B vssd1 vssd1 vccd1 vccd1 _5600_/A sky130_fd_sc_hd__nand2_2
X_7302_ _7398_/A _7303_/B vssd1 vssd1 vccd1 vccd1 _7327_/B sky130_fd_sc_hd__xnor2_1
X_4514_ _7908_/B _5617_/A vssd1 vssd1 vccd1 vccd1 _4541_/C sky130_fd_sc_hd__or2b_1
X_8282_ _8280_/A _8361_/A _8289_/B _8281_/Y vssd1 vssd1 vccd1 vccd1 _8287_/A sky130_fd_sc_hd__a2bb2o_2
X_5494_ _5494_/A vssd1 vssd1 vccd1 vccd1 _5558_/A sky130_fd_sc_hd__clkinv_2
X_4445_ _4451_/A vssd1 vssd1 vccd1 vccd1 _4450_/A sky130_fd_sc_hd__clkbuf_2
X_7233_ _7307_/B _7307_/C _7307_/A vssd1 vssd1 vccd1 vccd1 _7308_/A sky130_fd_sc_hd__o21a_1
X_4376_ _4377_/A vssd1 vssd1 vccd1 vccd1 _4376_/Y sky130_fd_sc_hd__inv_2
X_7164_ _7163_/A _7163_/B _7163_/C vssd1 vssd1 vccd1 vccd1 _7169_/B sky130_fd_sc_hd__a21o_1
XFILLER_58_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6115_ _6323_/D _6043_/A _6112_/X _6114_/X _6110_/B vssd1 vssd1 vccd1 vccd1 _6117_/A
+ sky130_fd_sc_hd__o221a_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7095_ _7095_/A _7095_/B vssd1 vssd1 vccd1 vccd1 _7096_/B sky130_fd_sc_hd__nor2_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6046_ _6046_/A _6046_/B vssd1 vssd1 vccd1 vccd1 _6046_/Y sky130_fd_sc_hd__xnor2_2
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7997_ _8069_/A _8069_/B vssd1 vssd1 vccd1 vccd1 _8074_/A sky130_fd_sc_hd__xnor2_1
XFILLER_54_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6948_ _7024_/A _6948_/B vssd1 vssd1 vccd1 vccd1 _7025_/B sky130_fd_sc_hd__nor2_1
X_6879_ _6787_/A _6787_/B _6878_/Y vssd1 vssd1 vccd1 vccd1 _6892_/A sky130_fd_sc_hd__a21o_1
X_8618_ input3/X _8618_/D vssd1 vssd1 vccd1 vccd1 _8618_/Q sky130_fd_sc_hd__dfxtp_1
X_8549_ _8546_/X _8547_/Y _8548_/Y _8564_/A vssd1 vssd1 vccd1 vccd1 _8549_/X sky130_fd_sc_hd__a211o_1
XFILLER_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7920_ _7920_/A _7920_/B vssd1 vssd1 vccd1 vccd1 _7921_/B sky130_fd_sc_hd__and2_1
X_7851_ _7851_/A vssd1 vssd1 vccd1 vccd1 _7851_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6802_ _7060_/A _7246_/B _6801_/Y _6728_/A vssd1 vssd1 vccd1 vccd1 _6803_/B sky130_fd_sc_hd__o211a_1
XFILLER_51_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7782_ _8714_/Q _7783_/A vssd1 vssd1 vccd1 vccd1 _8060_/A sky130_fd_sc_hd__or2b_1
X_4994_ _4994_/A _4994_/B vssd1 vssd1 vccd1 vccd1 _4995_/A sky130_fd_sc_hd__or2_1
X_6733_ _6734_/A _6734_/B _6734_/C vssd1 vssd1 vccd1 vccd1 _6735_/A sky130_fd_sc_hd__a21oi_1
XFILLER_51_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6664_ _6664_/A _6664_/B vssd1 vssd1 vccd1 vccd1 _6674_/A sky130_fd_sc_hd__nand2_1
XFILLER_31_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8403_ _8403_/A _8403_/B vssd1 vssd1 vccd1 vccd1 _8417_/A sky130_fd_sc_hd__xor2_2
X_5615_ _5615_/A _7783_/A vssd1 vssd1 vccd1 vccd1 _5616_/B sky130_fd_sc_hd__or2_1
X_6595_ _7296_/A _6580_/B _6773_/A vssd1 vssd1 vccd1 vccd1 _6596_/B sky130_fd_sc_hd__o21a_1
X_8334_ _8334_/A _8334_/B vssd1 vssd1 vccd1 vccd1 _8410_/C sky130_fd_sc_hd__xnor2_1
XFILLER_3_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5546_ _5549_/A _7871_/A vssd1 vssd1 vccd1 vccd1 _5546_/X sky130_fd_sc_hd__or2_1
X_8265_ _8267_/A _8267_/B vssd1 vssd1 vccd1 vccd1 _8503_/A sky130_fd_sc_hd__xnor2_1
X_5477_ _5477_/A _5477_/B vssd1 vssd1 vccd1 vccd1 _5533_/B sky130_fd_sc_hd__xnor2_4
X_7216_ _6995_/B _7214_/X _7213_/X _7210_/X vssd1 vssd1 vccd1 vccd1 _7217_/B sky130_fd_sc_hd__o211a_1
X_4428_ _4432_/A vssd1 vssd1 vccd1 vccd1 _4428_/Y sky130_fd_sc_hd__inv_2
X_8196_ _8196_/A _8361_/A vssd1 vssd1 vccd1 vccd1 _8196_/X sky130_fd_sc_hd__or2_1
X_7147_ _7147_/A _7147_/B vssd1 vssd1 vccd1 vccd1 _7147_/Y sky130_fd_sc_hd__nand2_1
XFILLER_98_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4359_ _4365_/A vssd1 vssd1 vccd1 vccd1 _4364_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_59_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7078_ _7078_/A _7078_/B _7078_/C vssd1 vssd1 vccd1 vccd1 _7081_/A sky130_fd_sc_hd__nor3_2
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8813__91 vssd1 vssd1 vccd1 vccd1 _8813__91/HI _8922_/A sky130_fd_sc_hd__conb_1
X_6029_ _6075_/A _6030_/B vssd1 vssd1 vccd1 vccd1 _6317_/A sky130_fd_sc_hd__or2_1
XFILLER_81_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5400_ _5421_/B vssd1 vssd1 vccd1 vccd1 _5433_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6380_ _8681_/Q vssd1 vssd1 vccd1 vccd1 _6459_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_5331_ _8627_/Q _6475_/B _5324_/B _8629_/Q vssd1 vssd1 vccd1 vccd1 _5332_/B sky130_fd_sc_hd__a31o_1
X_8050_ _8050_/A _8060_/B vssd1 vssd1 vccd1 vccd1 _8196_/A sky130_fd_sc_hd__nand2_2
X_7001_ _7001_/A _6962_/B vssd1 vssd1 vccd1 vccd1 _7001_/X sky130_fd_sc_hd__or2b_1
X_5262_ _4507_/X _4850_/A _4871_/A vssd1 vssd1 vccd1 vccd1 _5263_/B sky130_fd_sc_hd__o21a_1
X_5193_ _5193_/A _5193_/B _5193_/C _5193_/D vssd1 vssd1 vccd1 vccd1 _5193_/Y sky130_fd_sc_hd__nor4_1
XFILLER_83_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7903_ _7911_/B vssd1 vssd1 vccd1 vccd1 _8056_/B sky130_fd_sc_hd__buf_2
X_8883_ _8883_/A _4404_/Y vssd1 vssd1 vccd1 vccd1 io_out[30] sky130_fd_sc_hd__ebufn_8
X_7834_ _8051_/A _7988_/A vssd1 vssd1 vccd1 vccd1 _7836_/B sky130_fd_sc_hd__nand2_1
X_7765_ _7962_/B vssd1 vssd1 vccd1 vccd1 _8205_/B sky130_fd_sc_hd__clkbuf_2
X_6716_ _7160_/B _6718_/S _6641_/X vssd1 vssd1 vccd1 vccd1 _7060_/B sky130_fd_sc_hd__o21ai_4
X_4977_ _5004_/C _4977_/B vssd1 vssd1 vccd1 vccd1 _4977_/X sky130_fd_sc_hd__or2_1
XFILLER_11_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7696_ _8720_/Q _8596_/Q vssd1 vssd1 vccd1 vccd1 _7722_/B sky130_fd_sc_hd__xnor2_2
X_6647_ _6647_/A _7239_/A vssd1 vssd1 vccd1 vccd1 _6730_/A sky130_fd_sc_hd__nor2_1
X_6578_ _6815_/C vssd1 vssd1 vccd1 vccd1 _6647_/A sky130_fd_sc_hd__clkbuf_2
X_8317_ _8317_/A _8317_/B vssd1 vssd1 vccd1 vccd1 _8319_/B sky130_fd_sc_hd__nor2_1
XFILLER_3_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5529_ _5533_/B vssd1 vssd1 vccd1 vccd1 _6009_/A sky130_fd_sc_hd__clkbuf_2
X_8248_ _8293_/A _8248_/B vssd1 vssd1 vccd1 vccd1 _8251_/A sky130_fd_sc_hd__xor2_1
X_8179_ _8179_/A _8179_/B vssd1 vssd1 vccd1 vccd1 _8180_/B sky130_fd_sc_hd__nand2_1
XFILLER_86_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4900_ _5159_/B _5074_/B vssd1 vssd1 vccd1 vccd1 _5118_/C sky130_fd_sc_hd__or2_1
X_5880_ _6034_/A _5881_/B vssd1 vssd1 vccd1 vccd1 _5882_/A sky130_fd_sc_hd__nor2_1
X_4831_ _4831_/A _4831_/B _4831_/C vssd1 vssd1 vccd1 vccd1 _4960_/A sky130_fd_sc_hd__or3_1
XFILLER_33_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7550_ _8723_/Q vssd1 vssd1 vccd1 vccd1 _8566_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4762_ _4762_/A vssd1 vssd1 vccd1 vccd1 _8606_/D sky130_fd_sc_hd__clkbuf_1
X_7481_ _7480_/B _7480_/C _7480_/A vssd1 vssd1 vccd1 vccd1 _7481_/Y sky130_fd_sc_hd__a21oi_1
X_4693_ _4952_/A _4699_/B vssd1 vssd1 vccd1 vccd1 _4694_/A sky130_fd_sc_hd__or2_1
X_6501_ _8693_/Q vssd1 vssd1 vccd1 vccd1 _6539_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6432_ _6436_/C _6432_/B vssd1 vssd1 vccd1 vccd1 _8672_/D sky130_fd_sc_hd__nor2_1
X_8102_ _8088_/A _8088_/B _8101_/X vssd1 vssd1 vccd1 vccd1 _8186_/A sky130_fd_sc_hd__a21oi_1
X_6363_ _6375_/A _6371_/B vssd1 vssd1 vccd1 vccd1 _6367_/A sky130_fd_sc_hd__nor2_1
X_5314_ _8624_/Q _7533_/B vssd1 vssd1 vccd1 vccd1 _8624_/D sky130_fd_sc_hd__nor2_1
X_6294_ _6294_/A _6294_/B vssd1 vssd1 vccd1 vccd1 _6295_/B sky130_fd_sc_hd__xnor2_1
XFILLER_88_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8033_ _8117_/S vssd1 vssd1 vccd1 vccd1 _8317_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_5245_ _5245_/A _5245_/B _5245_/C _5245_/D vssd1 vssd1 vccd1 vccd1 _5245_/X sky130_fd_sc_hd__or4_1
XFILLER_102_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5176_ _5176_/A _5176_/B _5176_/C _5176_/D vssd1 vssd1 vccd1 vccd1 _5176_/X sky130_fd_sc_hd__or4_1
XFILLER_56_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8866_ _8866_/A _4382_/Y vssd1 vssd1 vccd1 vccd1 io_out[13] sky130_fd_sc_hd__ebufn_8
XFILLER_36_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7817_ _7904_/A vssd1 vssd1 vccd1 vccd1 _7817_/X sky130_fd_sc_hd__buf_2
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7748_ _7740_/A _7740_/B _7747_/X vssd1 vssd1 vccd1 vccd1 _7752_/B sky130_fd_sc_hd__a21oi_1
X_7679_ _7679_/A _7679_/B vssd1 vssd1 vccd1 vccd1 _7789_/B sky130_fd_sc_hd__and2_2
XFILLER_20_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5030_ _5235_/A _5174_/B _5030_/C _5219_/D vssd1 vssd1 vccd1 vccd1 _5030_/X sky130_fd_sc_hd__or4_1
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6981_ _7013_/A _7013_/B vssd1 vssd1 vccd1 vccd1 _6982_/B sky130_fd_sc_hd__xnor2_1
XFILLER_80_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8720_ input3/X _8720_/D vssd1 vssd1 vccd1 vccd1 _8720_/Q sky130_fd_sc_hd__dfxtp_1
X_5932_ _5932_/A _5932_/B vssd1 vssd1 vccd1 vccd1 _5933_/B sky130_fd_sc_hd__nand2_1
XFILLER_25_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5863_ _6072_/A _6072_/B vssd1 vssd1 vccd1 vccd1 _6074_/B sky130_fd_sc_hd__nor2_1
X_8651_ input3/X _8651_/D vssd1 vssd1 vccd1 vccd1 _8651_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7602_ _7603_/A _7603_/B vssd1 vssd1 vccd1 vccd1 _7602_/X sky130_fd_sc_hd__and2_1
X_4814_ _5115_/B vssd1 vssd1 vccd1 vccd1 _5153_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_8582_ input3/X _8582_/D vssd1 vssd1 vccd1 vccd1 _8582_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5794_ _5794_/A _5794_/B _5794_/C vssd1 vssd1 vccd1 vccd1 _5895_/B sky130_fd_sc_hd__and3_2
X_7533_ _7533_/A _7533_/B vssd1 vssd1 vccd1 vccd1 _7533_/Y sky130_fd_sc_hd__nor2_1
X_4745_ _4745_/A _5275_/B vssd1 vssd1 vccd1 vccd1 _4745_/Y sky130_fd_sc_hd__nand2_1
X_7464_ _7467_/A _7467_/B vssd1 vssd1 vccd1 vccd1 _7488_/B sky130_fd_sc_hd__xnor2_1
X_4676_ _4712_/B vssd1 vssd1 vccd1 vccd1 _4717_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7395_ _7395_/A _7395_/B _7395_/C vssd1 vssd1 vccd1 vccd1 _7480_/B sky130_fd_sc_hd__or3_2
X_6415_ _8668_/Q _6416_/B vssd1 vssd1 vccd1 vccd1 _6422_/C sky130_fd_sc_hd__and2_1
X_6346_ _6346_/A _8645_/Q vssd1 vssd1 vccd1 vccd1 _6347_/B sky130_fd_sc_hd__or2b_1
XFILLER_103_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8016_ _8093_/C vssd1 vssd1 vccd1 vccd1 _8499_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6277_ _6277_/A _6277_/B vssd1 vssd1 vccd1 vccd1 _6278_/B sky130_fd_sc_hd__xnor2_1
XFILLER_102_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5228_ _5075_/B _5227_/Y _4866_/A _5163_/B vssd1 vssd1 vccd1 vccd1 _5229_/C sky130_fd_sc_hd__a31o_1
XFILLER_29_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5159_ _5159_/A _5159_/B _5159_/C _5159_/D vssd1 vssd1 vccd1 vccd1 _5159_/X sky130_fd_sc_hd__or4_1
XFILLER_56_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8918_ _8918_/A _4443_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[27] sky130_fd_sc_hd__ebufn_8
X_8849_ _8849_/A _4362_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[28] sky130_fd_sc_hd__ebufn_8
XFILLER_72_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8774__52 vssd1 vssd1 vccd1 vccd1 _8774__52/HI _8883_/A sky130_fd_sc_hd__conb_1
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4530_ _5214_/A vssd1 vssd1 vccd1 vccd1 _5253_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_7_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4461_ _8599_/Q vssd1 vssd1 vccd1 vccd1 _7689_/B sky130_fd_sc_hd__inv_2
X_7180_ _7180_/A _7313_/A vssd1 vssd1 vccd1 vccd1 _7182_/B sky130_fd_sc_hd__xnor2_1
X_6200_ _6198_/Y _6023_/B _6199_/Y vssd1 vssd1 vccd1 vccd1 _6238_/A sky130_fd_sc_hd__a21bo_1
X_4392_ _4395_/A vssd1 vssd1 vccd1 vccd1 _4392_/Y sky130_fd_sc_hd__inv_2
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6131_ _6131_/A _6131_/B vssd1 vssd1 vccd1 vccd1 _6142_/B sky130_fd_sc_hd__xor2_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6062_ _6062_/A _6066_/B vssd1 vssd1 vccd1 vccd1 _6097_/A sky130_fd_sc_hd__xnor2_2
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5013_ _5068_/A _5118_/B _5215_/C vssd1 vssd1 vccd1 vccd1 _5014_/D sky130_fd_sc_hd__or3_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6964_ _6964_/A _6964_/B _6964_/C vssd1 vssd1 vccd1 vccd1 _6964_/Y sky130_fd_sc_hd__nor3_1
XFILLER_81_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6895_ _6895_/A _6852_/B vssd1 vssd1 vccd1 vccd1 _6895_/X sky130_fd_sc_hd__or2b_1
X_5915_ _5915_/A _5915_/B vssd1 vssd1 vccd1 vccd1 _5916_/B sky130_fd_sc_hd__xor2_1
X_8703_ input3/X _8703_/D vssd1 vssd1 vccd1 vccd1 _8703_/Q sky130_fd_sc_hd__dfxtp_1
X_8634_ input3/X _8634_/D vssd1 vssd1 vccd1 vccd1 _8634_/Q sky130_fd_sc_hd__dfxtp_1
X_5846_ _5753_/A _5751_/X _6180_/B _5674_/A vssd1 vssd1 vccd1 vccd1 _5921_/B sky130_fd_sc_hd__o22ai_2
XFILLER_21_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8565_ _8561_/A _7581_/X _8564_/Y _7541_/X vssd1 vssd1 vccd1 vccd1 _8724_/D sky130_fd_sc_hd__a211o_1
X_5777_ _5777_/A _5777_/B _5777_/C vssd1 vssd1 vccd1 vccd1 _5937_/A sky130_fd_sc_hd__and3_1
X_8496_ _8503_/B _8503_/C _8503_/A vssd1 vssd1 vccd1 vccd1 _8497_/C sky130_fd_sc_hd__a21oi_1
X_7516_ _8699_/Q _7516_/B vssd1 vssd1 vccd1 vccd1 _7516_/Y sky130_fd_sc_hd__xnor2_1
X_4728_ _4728_/A _4728_/B vssd1 vssd1 vccd1 vccd1 _5234_/A sky130_fd_sc_hd__nand2_1
X_7447_ _7470_/B _7470_/A vssd1 vssd1 vccd1 vccd1 _7447_/X sky130_fd_sc_hd__and2b_1
X_4659_ _4810_/A _4842_/C _4787_/B vssd1 vssd1 vccd1 vccd1 _4930_/A sky130_fd_sc_hd__or3_4
XFILLER_89_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7378_ _6647_/A _7378_/B _7418_/C _7378_/D vssd1 vssd1 vccd1 vccd1 _7385_/B sky130_fd_sc_hd__and4b_2
XFILLER_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6329_ _6341_/A _6301_/X _6326_/X _6328_/Y _6536_/B vssd1 vssd1 vccd1 vccd1 _6329_/X
+ sky130_fd_sc_hd__o41a_1
XFILLER_57_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5700_ _5980_/A vssd1 vssd1 vccd1 vccd1 _5956_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_16_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6680_ _6798_/B _7297_/B _7048_/C vssd1 vssd1 vccd1 vccd1 _6724_/B sky130_fd_sc_hd__or3_1
X_5631_ _5642_/A _5631_/B vssd1 vssd1 vccd1 vccd1 _5647_/A sky130_fd_sc_hd__nand2_2
X_8350_ _8429_/A _8429_/B vssd1 vssd1 vccd1 vccd1 _8427_/A sky130_fd_sc_hd__nand2_1
X_5562_ _5800_/A _6005_/B vssd1 vssd1 vccd1 vccd1 _5595_/B sky130_fd_sc_hd__nor2_1
X_8281_ _8306_/A vssd1 vssd1 vccd1 vccd1 _8281_/Y sky130_fd_sc_hd__inv_2
X_7301_ _7301_/A _7301_/B vssd1 vssd1 vccd1 vccd1 _7303_/B sky130_fd_sc_hd__xor2_1
X_4513_ _4782_/A _4513_/B vssd1 vssd1 vccd1 vccd1 _4542_/A sky130_fd_sc_hd__nor2_1
X_7232_ _7305_/A _7196_/X _7234_/A vssd1 vssd1 vccd1 vccd1 _7307_/A sky130_fd_sc_hd__o21ba_1
X_5493_ _5801_/C _5531_/B vssd1 vssd1 vccd1 vccd1 _5513_/A sky130_fd_sc_hd__xnor2_1
X_4444_ _4444_/A vssd1 vssd1 vccd1 vccd1 _4444_/Y sky130_fd_sc_hd__inv_2
X_4375_ _4377_/A vssd1 vssd1 vccd1 vccd1 _4375_/Y sky130_fd_sc_hd__inv_2
X_7163_ _7163_/A _7163_/B _7163_/C vssd1 vssd1 vccd1 vccd1 _7169_/A sky130_fd_sc_hd__nand3_1
X_7094_ _7088_/B _7114_/B _7092_/X _7306_/A vssd1 vssd1 vccd1 vccd1 _7096_/A sky130_fd_sc_hd__o22a_1
X_6114_ _6125_/A _6125_/B vssd1 vssd1 vccd1 vccd1 _6114_/X sky130_fd_sc_hd__and2_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6045_ _6323_/D _5755_/B _6043_/A vssd1 vssd1 vccd1 vccd1 _6109_/B sky130_fd_sc_hd__a21oi_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7996_ _7996_/A _7996_/B vssd1 vssd1 vccd1 vccd1 _8069_/B sky130_fd_sc_hd__xnor2_1
X_6947_ _6947_/A _6947_/B vssd1 vssd1 vccd1 vccd1 _6948_/B sky130_fd_sc_hd__and2_1
X_6878_ _6878_/A _6878_/B vssd1 vssd1 vccd1 vccd1 _6878_/Y sky130_fd_sc_hd__nor2_1
X_8617_ input3/X _8617_/D vssd1 vssd1 vccd1 vccd1 _8617_/Q sky130_fd_sc_hd__dfxtp_1
X_5829_ _5956_/A _5983_/A _5828_/B vssd1 vssd1 vccd1 vccd1 _5829_/Y sky130_fd_sc_hd__o21ai_1
X_8548_ _8546_/X _8547_/Y _6536_/B vssd1 vssd1 vccd1 vccd1 _8548_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_5_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8479_ _8479_/A _8479_/B vssd1 vssd1 vccd1 vccd1 _8480_/B sky130_fd_sc_hd__xnor2_1
XFILLER_78_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8744__22 vssd1 vssd1 vccd1 vccd1 _8744__22/HI _8839_/A sky130_fd_sc_hd__conb_1
XFILLER_32_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7850_ _7850_/A _7850_/B vssd1 vssd1 vccd1 vccd1 _7850_/X sky130_fd_sc_hd__or2_1
X_6801_ _6801_/A vssd1 vssd1 vccd1 vccd1 _6801_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7781_ _8050_/A _7671_/A _7796_/B _7685_/A vssd1 vssd1 vccd1 vccd1 _7902_/A sky130_fd_sc_hd__a31oi_4
XFILLER_51_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4993_ _5219_/D _4993_/B _4993_/C vssd1 vssd1 vccd1 vccd1 _4993_/X sky130_fd_sc_hd__or3_1
X_6732_ _6790_/A _6790_/B vssd1 vssd1 vccd1 vccd1 _6734_/C sky130_fd_sc_hd__xnor2_1
XFILLER_16_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6663_ _6671_/B vssd1 vssd1 vccd1 vccd1 _7177_/A sky130_fd_sc_hd__buf_2
XFILLER_31_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8402_ _8321_/A _8321_/B _8320_/A vssd1 vssd1 vccd1 vccd1 _8403_/B sky130_fd_sc_hd__a21oi_2
X_5614_ _5615_/A _7908_/B vssd1 vssd1 vccd1 vccd1 _5759_/A sky130_fd_sc_hd__nand2_2
X_6594_ _7226_/A _7236_/A vssd1 vssd1 vccd1 vccd1 _6773_/A sky130_fd_sc_hd__nor2_2
X_8333_ _8393_/B _8333_/B vssd1 vssd1 vccd1 vccd1 _8404_/A sky130_fd_sc_hd__xnor2_1
X_5545_ _5794_/A _5559_/B vssd1 vssd1 vccd1 vccd1 _6119_/A sky130_fd_sc_hd__nand2_2
X_8264_ _8264_/A _8264_/B vssd1 vssd1 vccd1 vccd1 _8267_/B sky130_fd_sc_hd__xnor2_1
XFILLER_2_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5476_ _5475_/A _5475_/B _5463_/A vssd1 vssd1 vccd1 vccd1 _5477_/A sky130_fd_sc_hd__a21o_1
X_7215_ _7210_/X _7213_/X _7214_/X _6995_/B vssd1 vssd1 vccd1 vccd1 _7217_/A sky130_fd_sc_hd__a211oi_1
X_8195_ _8383_/A vssd1 vssd1 vccd1 vccd1 _8385_/A sky130_fd_sc_hd__inv_2
X_4427_ _4427_/A vssd1 vssd1 vccd1 vccd1 _4432_/A sky130_fd_sc_hd__clkbuf_2
X_7146_ _7146_/A _7146_/B vssd1 vssd1 vccd1 vccd1 _7157_/A sky130_fd_sc_hd__xnor2_4
XFILLER_98_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4358_ _4358_/A vssd1 vssd1 vccd1 vccd1 _4358_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7077_ _7095_/B _7075_/X _7043_/Y _7044_/X vssd1 vssd1 vccd1 vccd1 _7078_/C sky130_fd_sc_hd__o211a_1
XFILLER_58_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6028_ _6170_/A _6028_/B vssd1 vssd1 vccd1 vccd1 _6030_/B sky130_fd_sc_hd__xnor2_1
XFILLER_46_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7979_ _8022_/B _7978_/C _7978_/A vssd1 vssd1 vccd1 vccd1 _7980_/C sky130_fd_sc_hd__a21o_1
XFILLER_54_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5330_ _8629_/Q _8628_/Q _5330_/C vssd1 vssd1 vccd1 vccd1 _5337_/C sky130_fd_sc_hd__and3_1
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5261_ _5261_/A _5261_/B _5261_/C _5260_/X vssd1 vssd1 vccd1 vccd1 _5269_/A sky130_fd_sc_hd__or4b_1
X_7000_ _7205_/A _6985_/B _6999_/X vssd1 vssd1 vccd1 vccd1 _7018_/A sky130_fd_sc_hd__o21ai_2
X_5192_ _5192_/A _5192_/B vssd1 vssd1 vccd1 vccd1 _5192_/Y sky130_fd_sc_hd__nor2_1
XFILLER_95_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7902_ _7902_/A _7902_/B vssd1 vssd1 vccd1 vccd1 _7998_/A sky130_fd_sc_hd__nor2_1
X_8882_ _8882_/A _4401_/Y vssd1 vssd1 vccd1 vccd1 io_out[29] sky130_fd_sc_hd__ebufn_8
XFILLER_36_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7833_ _7833_/A _7833_/B vssd1 vssd1 vccd1 vccd1 _7848_/A sky130_fd_sc_hd__xnor2_1
X_7764_ _7764_/A vssd1 vssd1 vccd1 vccd1 _7962_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_24_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6715_ _7020_/A _6978_/A vssd1 vssd1 vccd1 vccd1 _6951_/A sky130_fd_sc_hd__xnor2_2
X_4976_ _5174_/B _4976_/B _4976_/C _5054_/D vssd1 vssd1 vccd1 vccd1 _4977_/B sky130_fd_sc_hd__or4_1
X_7695_ _7695_/A vssd1 vssd1 vccd1 vccd1 _7722_/A sky130_fd_sc_hd__clkbuf_2
X_6646_ _7020_/A vssd1 vssd1 vccd1 vccd1 _7239_/A sky130_fd_sc_hd__buf_2
X_6577_ _7165_/A _7418_/B vssd1 vssd1 vccd1 vccd1 _6815_/C sky130_fd_sc_hd__nand2_1
X_8316_ _8224_/A _8224_/B _8315_/Y vssd1 vssd1 vccd1 vccd1 _8322_/A sky130_fd_sc_hd__o21ai_1
X_5528_ _5881_/B vssd1 vssd1 vccd1 vccd1 _5993_/A sky130_fd_sc_hd__buf_2
XFILLER_3_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8247_ _8292_/A _8292_/B vssd1 vssd1 vccd1 vccd1 _8248_/B sky130_fd_sc_hd__xor2_1
XFILLER_59_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5459_ _6375_/A _6777_/B vssd1 vssd1 vccd1 vccd1 _5460_/B sky130_fd_sc_hd__nor2_2
X_8178_ _8178_/A _8178_/B vssd1 vssd1 vccd1 vccd1 _8179_/B sky130_fd_sc_hd__or2_1
X_7129_ _7037_/A _7129_/B vssd1 vssd1 vccd1 vccd1 _7129_/X sky130_fd_sc_hd__and2b_1
XFILLER_74_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4830_ _5227_/A _4825_/Y _5109_/B _4829_/Y vssd1 vssd1 vccd1 vccd1 _5248_/A sky130_fd_sc_hd__a211o_2
XFILLER_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4761_ _5296_/A _4761_/B _4765_/B vssd1 vssd1 vccd1 vccd1 _4762_/A sky130_fd_sc_hd__and3_1
X_7480_ _7480_/A _7480_/B _7480_/C vssd1 vssd1 vccd1 vccd1 _7480_/X sky130_fd_sc_hd__and3_1
X_4692_ _4727_/A _5057_/A vssd1 vssd1 vccd1 vccd1 _4952_/A sky130_fd_sc_hd__nor2_1
X_6500_ _6536_/A _6505_/A _6497_/X _6531_/B vssd1 vssd1 vccd1 vccd1 _6500_/X sky130_fd_sc_hd__o31a_1
X_6431_ _8672_/Q _6429_/A _6409_/B vssd1 vssd1 vccd1 vccd1 _6432_/B sky130_fd_sc_hd__o21ai_1
X_6362_ _8661_/Q _5419_/X _6361_/Y _4743_/X vssd1 vssd1 vccd1 vccd1 _8661_/D sky130_fd_sc_hd__o211a_1
X_8101_ _8073_/A _8101_/B vssd1 vssd1 vccd1 vccd1 _8101_/X sky130_fd_sc_hd__and2b_1
X_5313_ _6511_/A vssd1 vssd1 vccd1 vccd1 _7533_/B sky130_fd_sc_hd__clkinv_2
X_6293_ _6197_/A _6197_/B _6292_/X vssd1 vssd1 vccd1 vccd1 _6294_/B sky130_fd_sc_hd__a21oi_1
X_8032_ _8107_/A _8107_/B vssd1 vssd1 vccd1 vccd1 _8041_/A sky130_fd_sc_hd__xnor2_1
XFILLER_88_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5244_ _5066_/A _5053_/D _5238_/X _5243_/X vssd1 vssd1 vccd1 vccd1 _5244_/X sky130_fd_sc_hd__o31a_1
X_5175_ _5175_/A _5175_/B vssd1 vssd1 vccd1 vccd1 _5176_/D sky130_fd_sc_hd__nand2_1
XFILLER_96_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8865_ _8865_/A _4381_/Y vssd1 vssd1 vccd1 vccd1 io_out[12] sky130_fd_sc_hd__ebufn_8
XFILLER_43_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7816_ _7816_/A _7816_/B vssd1 vssd1 vccd1 vccd1 _7833_/A sky130_fd_sc_hd__nand2_1
XFILLER_101_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7747_ _7747_/A _7747_/B vssd1 vssd1 vccd1 vccd1 _7747_/X sky130_fd_sc_hd__or2_1
X_4959_ _4959_/A vssd1 vssd1 vccd1 vccd1 _5145_/B sky130_fd_sc_hd__buf_2
XFILLER_24_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7678_ _7643_/A _7643_/B _7641_/B _7657_/X _7639_/X vssd1 vssd1 vccd1 vccd1 _7679_/B
+ sky130_fd_sc_hd__a311o_1
XFILLER_20_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6629_ _6629_/A vssd1 vssd1 vccd1 vccd1 _6798_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_10_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6980_ _6980_/A _6980_/B vssd1 vssd1 vccd1 vccd1 _7013_/B sky130_fd_sc_hd__xnor2_1
X_5931_ _5932_/A _5932_/B vssd1 vssd1 vccd1 vccd1 _5976_/A sky130_fd_sc_hd__nor2_1
XFILLER_25_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8650_ input3/X _8650_/D vssd1 vssd1 vccd1 vccd1 _8650_/Q sky130_fd_sc_hd__dfxtp_1
X_5862_ _5862_/A _5862_/B vssd1 vssd1 vccd1 vccd1 _6072_/B sky130_fd_sc_hd__xnor2_1
X_7601_ _7594_/A _7596_/B _7594_/B vssd1 vssd1 vccd1 vccd1 _7603_/B sky130_fd_sc_hd__o21ba_1
X_4813_ _5172_/B vssd1 vssd1 vccd1 vccd1 _5115_/B sky130_fd_sc_hd__clkbuf_2
X_8581_ input3/X _8581_/D vssd1 vssd1 vccd1 vccd1 _8581_/Q sky130_fd_sc_hd__dfxtp_1
X_5793_ _5997_/A _5729_/B _5792_/X vssd1 vssd1 vccd1 vccd1 _5889_/B sky130_fd_sc_hd__a21oi_2
X_4744_ _4850_/B _4733_/Y _5275_/B _4824_/C _4743_/X vssd1 vssd1 vccd1 vccd1 _8603_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_21_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7532_ _7532_/A _7532_/B vssd1 vssd1 vccd1 vccd1 _7532_/X sky130_fd_sc_hd__or2_1
X_7463_ _7462_/A _7218_/B _7217_/A vssd1 vssd1 vccd1 vccd1 _7467_/B sky130_fd_sc_hd__a21o_1
X_4675_ _6507_/A _4675_/B vssd1 vssd1 vccd1 vccd1 _4712_/B sky130_fd_sc_hd__nor2_1
X_7394_ _7396_/A _7396_/B vssd1 vssd1 vccd1 vccd1 _7395_/C sky130_fd_sc_hd__and2_1
X_6414_ _6414_/A vssd1 vssd1 vccd1 vccd1 _8667_/D sky130_fd_sc_hd__clkbuf_1
X_6345_ _8645_/Q _6346_/A vssd1 vssd1 vccd1 vccd1 _6347_/A sky130_fd_sc_hd__or2b_1
X_6276_ _6238_/A _6238_/B _6275_/X vssd1 vssd1 vccd1 vccd1 _6278_/A sky130_fd_sc_hd__a21oi_1
X_8015_ _8015_/A _8015_/B _8015_/C vssd1 vssd1 vccd1 vccd1 _8093_/C sky130_fd_sc_hd__nand3_1
X_5227_ _5227_/A _5227_/B vssd1 vssd1 vccd1 vccd1 _5227_/Y sky130_fd_sc_hd__nand2_1
XFILLER_102_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5158_ _5092_/C _5153_/B _5156_/Y _5157_/Y vssd1 vssd1 vccd1 vccd1 _5159_/D sky130_fd_sc_hd__o31a_1
XFILLER_29_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5089_ _5229_/D _5230_/A vssd1 vssd1 vccd1 vccd1 _5089_/Y sky130_fd_sc_hd__nand2_1
X_8917_ _8917_/A _4442_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[26] sky130_fd_sc_hd__ebufn_8
XFILLER_56_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8848_ _8848_/A _4361_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[27] sky130_fd_sc_hd__ebufn_8
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4460_ _8600_/Q vssd1 vssd1 vccd1 vccd1 _7753_/A sky130_fd_sc_hd__buf_2
XFILLER_7_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4391_ _4395_/A vssd1 vssd1 vccd1 vccd1 _4391_/Y sky130_fd_sc_hd__clkinv_2
X_6130_ _6131_/A _6131_/B vssd1 vssd1 vccd1 vccd1 _6140_/B sky130_fd_sc_hd__nor2_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6061_ _6061_/A _6061_/B vssd1 vssd1 vccd1 vccd1 _6066_/B sky130_fd_sc_hd__xor2_2
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5012_ _5012_/A vssd1 vssd1 vccd1 vccd1 _5215_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_38_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6963_ _6963_/A _6963_/B vssd1 vssd1 vccd1 vccd1 _6964_/C sky130_fd_sc_hd__xnor2_1
XFILLER_53_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6894_ _7159_/A _7159_/B vssd1 vssd1 vccd1 vccd1 _6894_/Y sky130_fd_sc_hd__nor2_1
XFILLER_81_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8702_ input3/X _8702_/D vssd1 vssd1 vccd1 vccd1 _8702_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5914_ _5914_/A _5914_/B vssd1 vssd1 vccd1 vccd1 _5915_/B sky130_fd_sc_hd__xor2_1
X_8633_ input3/X _8633_/D vssd1 vssd1 vccd1 vccd1 _8633_/Q sky130_fd_sc_hd__dfxtp_1
X_5845_ _5845_/A _5865_/B vssd1 vssd1 vccd1 vccd1 _5859_/A sky130_fd_sc_hd__xnor2_1
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8564_ _8564_/A _8564_/B vssd1 vssd1 vccd1 vccd1 _8564_/Y sky130_fd_sc_hd__nor2_1
X_5776_ _5675_/B _5755_/B _5983_/A vssd1 vssd1 vccd1 vccd1 _5777_/C sky130_fd_sc_hd__o21a_1
X_8495_ _8495_/A vssd1 vssd1 vccd1 vccd1 _8497_/A sky130_fd_sc_hd__inv_2
X_7515_ _7515_/A _7515_/B vssd1 vssd1 vccd1 vccd1 _7516_/B sky130_fd_sc_hd__nand2_1
XFILLER_21_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4727_ _4727_/A vssd1 vssd1 vccd1 vccd1 _4728_/A sky130_fd_sc_hd__clkbuf_2
X_7446_ _7446_/A _7446_/B vssd1 vssd1 vccd1 vccd1 _7470_/A sky130_fd_sc_hd__xnor2_1
X_4658_ _5607_/B _4831_/B vssd1 vssd1 vccd1 vccd1 _4787_/B sky130_fd_sc_hd__nand2_1
X_7377_ _7377_/A _7377_/B vssd1 vssd1 vccd1 vccd1 _7385_/A sky130_fd_sc_hd__xor2_1
XFILLER_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4589_ _8572_/Q _8571_/Q _8573_/Q vssd1 vssd1 vccd1 vccd1 _4598_/C sky130_fd_sc_hd__and3_1
XFILLER_88_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6328_ _6302_/A _6332_/B _6304_/X vssd1 vssd1 vccd1 vccd1 _6328_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_103_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6259_ _6259_/A _6259_/B vssd1 vssd1 vccd1 vccd1 _6260_/B sky130_fd_sc_hd__xnor2_1
XFILLER_76_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5630_ _5646_/A vssd1 vssd1 vccd1 vccd1 _5826_/A sky130_fd_sc_hd__clkbuf_2
X_5561_ _5561_/A vssd1 vssd1 vccd1 vccd1 _6005_/B sky130_fd_sc_hd__clkbuf_2
X_8280_ _8280_/A _8306_/B vssd1 vssd1 vccd1 vccd1 _8289_/B sky130_fd_sc_hd__xor2_1
X_7300_ _7300_/A _7315_/C vssd1 vssd1 vccd1 vccd1 _7301_/B sky130_fd_sc_hd__xnor2_1
X_5492_ _5512_/A _5492_/B vssd1 vssd1 vccd1 vccd1 _5531_/B sky130_fd_sc_hd__xnor2_1
X_4512_ _4495_/A _4518_/C _4495_/B _4781_/A vssd1 vssd1 vccd1 vccd1 _4513_/B sky130_fd_sc_hd__o211a_1
X_7231_ _7231_/A _7376_/A _7230_/X vssd1 vssd1 vccd1 vccd1 _7307_/C sky130_fd_sc_hd__nor3b_1
XFILLER_7_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4443_ _4444_/A vssd1 vssd1 vccd1 vccd1 _4443_/Y sky130_fd_sc_hd__inv_2
X_4374_ _4377_/A vssd1 vssd1 vccd1 vccd1 _4374_/Y sky130_fd_sc_hd__inv_2
X_7162_ _7266_/A _7162_/B vssd1 vssd1 vccd1 vccd1 _7262_/A sky130_fd_sc_hd__xor2_1
XFILLER_98_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7093_ _7220_/A vssd1 vssd1 vccd1 vccd1 _7306_/A sky130_fd_sc_hd__clkinv_2
X_6113_ _6123_/B _6113_/B vssd1 vssd1 vccd1 vccd1 _6125_/B sky130_fd_sc_hd__xnor2_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6044_ _6044_/A _6044_/B _5749_/B vssd1 vssd1 vccd1 vccd1 _6108_/A sky130_fd_sc_hd__or3b_2
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7995_ _8057_/A _7995_/B vssd1 vssd1 vccd1 vccd1 _7996_/B sky130_fd_sc_hd__nor2_1
X_6946_ _6947_/A _6947_/B vssd1 vssd1 vccd1 vccd1 _7024_/A sky130_fd_sc_hd__nor2_1
XFILLER_54_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6877_ _7151_/A _7205_/B _6876_/X vssd1 vssd1 vccd1 vccd1 _6893_/A sky130_fd_sc_hd__a21bo_1
XFILLER_34_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8616_ input3/X _8616_/D vssd1 vssd1 vccd1 vccd1 _8616_/Q sky130_fd_sc_hd__dfxtp_1
X_5828_ _5828_/A _5828_/B vssd1 vssd1 vccd1 vccd1 _5831_/A sky130_fd_sc_hd__xnor2_1
X_8547_ _8542_/A _8542_/B _8540_/A vssd1 vssd1 vccd1 vccd1 _8547_/Y sky130_fd_sc_hd__a21oi_1
X_5759_ _5759_/A _5826_/A vssd1 vssd1 vccd1 vccd1 _6284_/S sky130_fd_sc_hd__nand2_2
X_8478_ _8375_/A _8476_/Y _8477_/X vssd1 vssd1 vccd1 vccd1 _8479_/B sky130_fd_sc_hd__a21oi_1
X_7429_ _7434_/A _7434_/B _7428_/X vssd1 vssd1 vccd1 vccd1 _7449_/C sky130_fd_sc_hd__o21ai_1
XFILLER_78_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6800_ _7048_/A _7048_/C vssd1 vssd1 vccd1 vccd1 _6801_/A sky130_fd_sc_hd__nor2_1
XFILLER_90_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7780_ _8283_/A _8305_/A vssd1 vssd1 vccd1 vccd1 _7796_/B sky130_fd_sc_hd__nor2_2
X_4992_ _5176_/A _5241_/A _5241_/B _5151_/B vssd1 vssd1 vccd1 vccd1 _4993_/C sky130_fd_sc_hd__or4_1
X_6731_ _6827_/A _6731_/B vssd1 vssd1 vccd1 vccd1 _6790_/B sky130_fd_sc_hd__xnor2_2
XFILLER_51_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6662_ _6687_/A _6687_/B vssd1 vssd1 vccd1 vccd1 _6671_/B sky130_fd_sc_hd__xnor2_1
X_8401_ _8401_/A _8401_/B vssd1 vssd1 vccd1 vccd1 _8403_/A sky130_fd_sc_hd__nand2_1
X_5613_ _6044_/A vssd1 vssd1 vccd1 vccd1 _6123_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_8332_ _8126_/B _8407_/S _8331_/Y _8222_/A vssd1 vssd1 vccd1 vccd1 _8333_/B sky130_fd_sc_hd__o2bb2a_1
X_6593_ _6593_/A vssd1 vssd1 vccd1 vccd1 _7226_/A sky130_fd_sc_hd__clkbuf_2
X_5544_ _5993_/A _6005_/A vssd1 vssd1 vccd1 vccd1 _5553_/A sky130_fd_sc_hd__nor2_1
X_8263_ _8263_/A _8263_/B vssd1 vssd1 vccd1 vccd1 _8267_/A sky130_fd_sc_hd__nand2_1
X_5475_ _5475_/A _5475_/B vssd1 vssd1 vccd1 vccd1 _5494_/A sky130_fd_sc_hd__xnor2_2
X_7214_ _6995_/A _6993_/Y _6991_/X _6992_/X vssd1 vssd1 vccd1 vccd1 _7214_/X sky130_fd_sc_hd__o211a_1
X_4426_ _4426_/A vssd1 vssd1 vccd1 vccd1 _4426_/Y sky130_fd_sc_hd__clkinv_4
X_8194_ _8194_/A _8194_/B vssd1 vssd1 vccd1 vccd1 _8201_/A sky130_fd_sc_hd__and2_1
X_7145_ _7145_/A _7145_/B vssd1 vssd1 vccd1 vccd1 _7146_/B sky130_fd_sc_hd__xnor2_2
X_4357_ _4358_/A vssd1 vssd1 vccd1 vccd1 _4357_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7076_ _7043_/Y _7044_/X _7095_/B _7075_/X vssd1 vssd1 vccd1 vccd1 _7078_/B sky130_fd_sc_hd__a211oi_4
XFILLER_58_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6027_ _6027_/A _6027_/B vssd1 vssd1 vccd1 vccd1 _6028_/B sky130_fd_sc_hd__xor2_1
XFILLER_39_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7978_ _7978_/A _8022_/B _7978_/C vssd1 vssd1 vccd1 vccd1 _8021_/A sky130_fd_sc_hd__nand3_1
X_6929_ _6977_/S vssd1 vssd1 vccd1 vccd1 _7065_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_10_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8804__82 vssd1 vssd1 vccd1 vccd1 _8804__82/HI _8913_/A sky130_fd_sc_hd__conb_1
XFILLER_64_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5260_ _5234_/X _5251_/X _5259_/X _5190_/A vssd1 vssd1 vccd1 vccd1 _5260_/X sky130_fd_sc_hd__a31o_1
XFILLER_68_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5191_ _5191_/A _5192_/B vssd1 vssd1 vccd1 vccd1 _5203_/A sky130_fd_sc_hd__nor2_1
XFILLER_95_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7901_ _7948_/B _7948_/C _7948_/A vssd1 vssd1 vccd1 vccd1 _7929_/B sky130_fd_sc_hd__a21o_1
XFILLER_55_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8881_ _8881_/A _4400_/Y vssd1 vssd1 vccd1 vccd1 io_out[28] sky130_fd_sc_hd__ebufn_8
XFILLER_70_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7832_ _7944_/A _7832_/B vssd1 vssd1 vccd1 vccd1 _7845_/A sky130_fd_sc_hd__xor2_1
X_7763_ _8229_/A vssd1 vssd1 vccd1 vccd1 _8331_/A sky130_fd_sc_hd__clkbuf_2
X_4975_ _8592_/Q _4975_/B vssd1 vssd1 vccd1 vccd1 _5054_/D sky130_fd_sc_hd__nand2_1
XFILLER_24_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6714_ _6806_/A _6806_/B vssd1 vssd1 vccd1 vccd1 _6978_/A sky130_fd_sc_hd__nor2_4
X_7694_ _8595_/Q _8719_/Q vssd1 vssd1 vccd1 vccd1 _7695_/A sky130_fd_sc_hd__or2b_1
X_6645_ _6645_/A _6718_/S vssd1 vssd1 vccd1 vccd1 _7065_/A sky130_fd_sc_hd__xnor2_2
X_6576_ _7176_/A vssd1 vssd1 vccd1 vccd1 _7418_/B sky130_fd_sc_hd__clkbuf_2
X_8315_ _8315_/A _8315_/B vssd1 vssd1 vccd1 vccd1 _8315_/Y sky130_fd_sc_hd__nand2_1
X_5527_ _6033_/A _6033_/B _5526_/X vssd1 vssd1 vccd1 vccd1 _5571_/A sky130_fd_sc_hd__a21o_1
X_8246_ _8147_/A _8384_/A _8146_/B _8151_/A _8151_/B vssd1 vssd1 vccd1 vccd1 _8292_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_78_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5458_ _8662_/Q vssd1 vssd1 vccd1 vccd1 _6375_/A sky130_fd_sc_hd__inv_2
X_8177_ _8178_/A _8178_/B vssd1 vssd1 vccd1 vccd1 _8179_/A sky130_fd_sc_hd__nand2_1
X_4409_ _4427_/A vssd1 vssd1 vccd1 vccd1 _4414_/A sky130_fd_sc_hd__clkbuf_2
X_5389_ _5549_/A _5402_/C _6371_/B vssd1 vssd1 vccd1 vccd1 _5389_/Y sky130_fd_sc_hd__o21ai_1
X_7128_ _7128_/A _7128_/B vssd1 vssd1 vccd1 vccd1 _7132_/A sky130_fd_sc_hd__xnor2_1
XFILLER_86_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7059_ _7058_/A _7058_/B _7058_/C vssd1 vssd1 vccd1 vccd1 _7074_/B sky130_fd_sc_hd__a21oi_1
XFILLER_74_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4760_ _4760_/A _4856_/A _4495_/A vssd1 vssd1 vccd1 vccd1 _4765_/B sky130_fd_sc_hd__or3b_1
XFILLER_81_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4691_ _5185_/A vssd1 vssd1 vccd1 vccd1 _5057_/A sky130_fd_sc_hd__clkbuf_2
X_6430_ _6430_/A _8672_/Q _6430_/C vssd1 vssd1 vccd1 vccd1 _6436_/C sky130_fd_sc_hd__and3_1
X_6361_ _6358_/X _6359_/Y _6360_/Y vssd1 vssd1 vccd1 vccd1 _6361_/Y sky130_fd_sc_hd__o21ai_1
X_8100_ _8090_/A _8090_/B _8099_/X vssd1 vssd1 vccd1 vccd1 _8264_/A sky130_fd_sc_hd__a21o_1
X_5312_ _5320_/A vssd1 vssd1 vccd1 vccd1 _6511_/A sky130_fd_sc_hd__clkbuf_2
X_6292_ _6194_/B _6292_/B vssd1 vssd1 vccd1 vccd1 _6292_/X sky130_fd_sc_hd__and2b_1
X_8031_ _8031_/A _8031_/B vssd1 vssd1 vccd1 vccd1 _8107_/B sky130_fd_sc_hd__xnor2_1
X_5243_ _5243_/A _5243_/B _5243_/C _5243_/D vssd1 vssd1 vccd1 vccd1 _5243_/X sky130_fd_sc_hd__or4_1
XFILLER_102_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5174_ _5240_/B _5174_/B vssd1 vssd1 vccd1 vccd1 _5175_/A sky130_fd_sc_hd__nor2_1
XFILLER_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8795__73 vssd1 vssd1 vccd1 vccd1 _8795__73/HI _8904_/A sky130_fd_sc_hd__conb_1
X_8864_ _8864_/A _4380_/Y vssd1 vssd1 vccd1 vccd1 io_out[11] sky130_fd_sc_hd__ebufn_8
X_7815_ _7815_/A _7815_/B vssd1 vssd1 vccd1 vccd1 _7829_/A sky130_fd_sc_hd__nand2_1
XFILLER_52_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7746_ _7746_/A _7864_/A vssd1 vssd1 vccd1 vccd1 _7757_/A sky130_fd_sc_hd__nand2_1
XFILLER_51_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4958_ _5166_/A vssd1 vssd1 vccd1 vccd1 _5219_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_24_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7677_ _7677_/A _7676_/X vssd1 vssd1 vccd1 vccd1 _7789_/A sky130_fd_sc_hd__or2b_4
X_4889_ _5143_/A vssd1 vssd1 vccd1 vccd1 _5231_/A sky130_fd_sc_hd__clkbuf_2
X_6628_ _6628_/A _7783_/A vssd1 vssd1 vccd1 vccd1 _6629_/A sky130_fd_sc_hd__and2_1
X_6559_ _6710_/A vssd1 vssd1 vccd1 vccd1 _6561_/A sky130_fd_sc_hd__inv_2
X_8229_ _8229_/A _8334_/B vssd1 vssd1 vccd1 vccd1 _8232_/A sky130_fd_sc_hd__xnor2_1
XFILLER_10_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5930_ _5777_/B _5852_/B _5850_/Y vssd1 vssd1 vccd1 vccd1 _5932_/B sky130_fd_sc_hd__a21o_1
XFILLER_18_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7600_ _7604_/A _7615_/B vssd1 vssd1 vccd1 vccd1 _7603_/A sky130_fd_sc_hd__xnor2_1
X_5861_ _5861_/A _5861_/B _5709_/C vssd1 vssd1 vccd1 vccd1 _6072_/A sky130_fd_sc_hd__or3b_1
X_4812_ _4839_/B _4897_/C vssd1 vssd1 vccd1 vccd1 _5172_/B sky130_fd_sc_hd__nor2_2
X_8580_ input3/X _8580_/D vssd1 vssd1 vccd1 vccd1 _8580_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5792_ _5792_/A _5792_/B vssd1 vssd1 vccd1 vccd1 _5792_/X sky130_fd_sc_hd__and2_1
X_7531_ _7532_/A _7532_/B vssd1 vssd1 vccd1 vccd1 _7543_/A sky130_fd_sc_hd__nand2_1
X_4743_ _5296_/A vssd1 vssd1 vccd1 vccd1 _4743_/X sky130_fd_sc_hd__buf_2
X_7462_ _7462_/A _7462_/B vssd1 vssd1 vccd1 vccd1 _7467_/A sky130_fd_sc_hd__xnor2_1
X_4674_ _4732_/A _4732_/B _5113_/A _4681_/B vssd1 vssd1 vccd1 vccd1 _4675_/B sky130_fd_sc_hd__and4bb_1
X_6413_ _6416_/B _6413_/B _6468_/B vssd1 vssd1 vccd1 vccd1 _6414_/A sky130_fd_sc_hd__and3b_1
X_7393_ _7393_/A _7393_/B vssd1 vssd1 vccd1 vccd1 _7396_/B sky130_fd_sc_hd__xor2_1
X_6344_ _6344_/A vssd1 vssd1 vccd1 vccd1 _8658_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6275_ _6239_/A _6275_/B vssd1 vssd1 vccd1 vccd1 _6275_/X sky130_fd_sc_hd__and2b_1
XFILLER_102_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8014_ _8017_/A _8013_/C _8013_/A vssd1 vssd1 vccd1 vccd1 _8015_/C sky130_fd_sc_hd__o21ai_1
X_5226_ _5226_/A _5226_/B vssd1 vssd1 vccd1 vccd1 _5261_/C sky130_fd_sc_hd__nand2_1
XFILLER_102_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5157_ _4930_/A _4930_/B _5152_/Y _5105_/A _5219_/A vssd1 vssd1 vccd1 vccd1 _5157_/Y
+ sky130_fd_sc_hd__o221ai_1
X_5088_ _5071_/A _5256_/A _5135_/C _4941_/C _5087_/X vssd1 vssd1 vccd1 vccd1 _5088_/X
+ sky130_fd_sc_hd__o32a_1
X_8916_ _8916_/A _4441_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[25] sky130_fd_sc_hd__ebufn_8
XFILLER_56_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8847_ _8847_/A _4360_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[26] sky130_fd_sc_hd__ebufn_8
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7729_ _7885_/A _7729_/B vssd1 vssd1 vccd1 vccd1 _7814_/B sky130_fd_sc_hd__xnor2_1
XFILLER_8_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4390_ _4396_/A vssd1 vssd1 vccd1 vccd1 _4395_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_7_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6060_ _6060_/A _6060_/B vssd1 vssd1 vccd1 vccd1 _6062_/A sky130_fd_sc_hd__nor2_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5011_ _5011_/A _5041_/B vssd1 vssd1 vccd1 vccd1 _5012_/A sky130_fd_sc_hd__nor2_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6962_ _7001_/A _6962_/B vssd1 vssd1 vccd1 vccd1 _6963_/B sky130_fd_sc_hd__xnor2_1
XFILLER_53_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8765__43 vssd1 vssd1 vccd1 vccd1 _8765__43/HI _8860_/A sky130_fd_sc_hd__conb_1
X_6893_ _6893_/A _6992_/A vssd1 vssd1 vccd1 vccd1 _7159_/B sky130_fd_sc_hd__xor2_1
X_8701_ input3/X _8701_/D vssd1 vssd1 vccd1 vccd1 _8701_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5913_ _5913_/A _5913_/B vssd1 vssd1 vccd1 vccd1 _5914_/B sky130_fd_sc_hd__nor2_1
X_8632_ input3/X _8632_/D vssd1 vssd1 vccd1 vccd1 _8632_/Q sky130_fd_sc_hd__dfxtp_1
X_5844_ _5844_/A _5844_/B vssd1 vssd1 vccd1 vccd1 _5865_/B sky130_fd_sc_hd__xor2_1
XFILLER_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8563_ _8563_/A _8563_/B vssd1 vssd1 vccd1 vccd1 _8564_/B sky130_fd_sc_hd__xnor2_1
X_7514_ _7514_/A _8686_/Q vssd1 vssd1 vccd1 vccd1 _7515_/B sky130_fd_sc_hd__or2b_1
X_5775_ _5826_/B vssd1 vssd1 vccd1 vccd1 _5983_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_21_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8494_ _8491_/Y _8492_/X _8493_/X vssd1 vssd1 vccd1 vccd1 _8494_/X sky130_fd_sc_hd__o21a_1
X_4726_ _4810_/B vssd1 vssd1 vccd1 vccd1 _4909_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7445_ _7494_/A _7495_/A _7495_/B _7442_/B _7442_/A vssd1 vssd1 vccd1 vccd1 _7470_/B
+ sky130_fd_sc_hd__o32a_1
X_4657_ _4657_/A vssd1 vssd1 vccd1 vccd1 _4661_/A sky130_fd_sc_hd__clkbuf_2
X_7376_ _7376_/A _7231_/A vssd1 vssd1 vccd1 vccd1 _7380_/A sky130_fd_sc_hd__or2b_1
XFILLER_1_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4588_ _4588_/A vssd1 vssd1 vccd1 vccd1 _8572_/D sky130_fd_sc_hd__clkbuf_1
X_6327_ _6327_/A _6327_/B vssd1 vssd1 vccd1 vccd1 _6332_/B sky130_fd_sc_hd__xor2_1
XFILLER_103_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6258_ _5993_/A _5551_/A _5549_/Y _5794_/B _5488_/Y vssd1 vssd1 vccd1 vccd1 _6259_/B
+ sky130_fd_sc_hd__o2111a_1
XFILLER_103_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6189_ _6189_/A _6189_/B vssd1 vssd1 vccd1 vccd1 _6192_/A sky130_fd_sc_hd__xnor2_1
X_5209_ _4953_/X _5179_/X _5190_/X _5208_/X _4707_/B vssd1 vssd1 vccd1 vccd1 _5209_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_72_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5560_ _5560_/A _5560_/B vssd1 vssd1 vccd1 vccd1 _5567_/B sky130_fd_sc_hd__and2_1
X_4511_ _5617_/A vssd1 vssd1 vccd1 vccd1 _4781_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5491_ _6213_/A _5539_/B _5488_/Y _6034_/B vssd1 vssd1 vccd1 vccd1 _5492_/B sky130_fd_sc_hd__o211a_1
X_4442_ _4444_/A vssd1 vssd1 vccd1 vccd1 _4442_/Y sky130_fd_sc_hd__inv_2
X_7230_ _7230_/A _7434_/A vssd1 vssd1 vccd1 vccd1 _7230_/X sky130_fd_sc_hd__xor2_1
XFILLER_104_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4373_ _4377_/A vssd1 vssd1 vccd1 vccd1 _4373_/Y sky130_fd_sc_hd__inv_2
X_7161_ _7161_/A _7161_/B vssd1 vssd1 vccd1 vccd1 _7162_/B sky130_fd_sc_hd__nor2_1
X_7092_ _7092_/A _7236_/B _7092_/C vssd1 vssd1 vccd1 vccd1 _7092_/X sky130_fd_sc_hd__or3_1
X_6112_ _6123_/B _6113_/B vssd1 vssd1 vccd1 vccd1 _6112_/X sky130_fd_sc_hd__and2b_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6043_ _6043_/A vssd1 vssd1 vccd1 vccd1 _6044_/B sky130_fd_sc_hd__inv_2
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7994_ _8068_/A _8068_/B vssd1 vssd1 vccd1 vccd1 _8069_/A sky130_fd_sc_hd__xnor2_1
X_6945_ _6804_/A _6804_/B _6803_/B _6944_/Y vssd1 vssd1 vccd1 vccd1 _7001_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_41_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6876_ _6876_/A _6876_/B _6876_/C vssd1 vssd1 vccd1 vccd1 _6876_/X sky130_fd_sc_hd__or3_1
XFILLER_34_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5827_ _5983_/B _5870_/B vssd1 vssd1 vccd1 vccd1 _5828_/B sky130_fd_sc_hd__xnor2_2
XFILLER_22_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8615_ input3/X _8615_/D vssd1 vssd1 vccd1 vccd1 _8615_/Q sky130_fd_sc_hd__dfxtp_1
X_8546_ _8546_/A _8561_/B vssd1 vssd1 vccd1 vccd1 _8546_/X sky130_fd_sc_hd__xor2_1
X_5758_ _5922_/A _6110_/B vssd1 vssd1 vccd1 vccd1 _5954_/B sky130_fd_sc_hd__nand2_1
XFILLER_22_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8477_ _8372_/B _8477_/B vssd1 vssd1 vccd1 vccd1 _8477_/X sky130_fd_sc_hd__and2b_1
X_4709_ _4709_/A _5113_/A vssd1 vssd1 vccd1 vccd1 _4786_/B sky130_fd_sc_hd__nand2_1
X_7428_ _7428_/A _7428_/B vssd1 vssd1 vccd1 vccd1 _7428_/X sky130_fd_sc_hd__or2_1
X_5689_ _6323_/C _5980_/A vssd1 vssd1 vccd1 vccd1 _6046_/A sky130_fd_sc_hd__nor2_1
X_7359_ _7368_/B _7368_/A vssd1 vssd1 vccd1 vccd1 _7366_/C sky130_fd_sc_hd__or2b_1
XFILLER_103_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6730_ _6730_/A _6730_/B vssd1 vssd1 vccd1 vccd1 _6731_/B sky130_fd_sc_hd__xnor2_1
XFILLER_51_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4991_ _5143_/B _5092_/C _5176_/B _4990_/Y _5092_/A vssd1 vssd1 vccd1 vccd1 _4993_/B
+ sky130_fd_sc_hd__o32a_1
XFILLER_90_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8735__13 vssd1 vssd1 vccd1 vccd1 _8735__13/HI _8830_/A sky130_fd_sc_hd__conb_1
X_6661_ _6581_/A _6581_/B _6620_/A vssd1 vssd1 vccd1 vccd1 _6687_/B sky130_fd_sc_hd__a21boi_1
X_8400_ _8400_/A _8400_/B _8400_/C vssd1 vssd1 vccd1 vccd1 _8401_/B sky130_fd_sc_hd__or3_1
X_6592_ _6592_/A _6592_/B vssd1 vssd1 vccd1 vccd1 _6593_/A sky130_fd_sc_hd__and2_1
X_5612_ _5671_/A vssd1 vssd1 vccd1 vccd1 _6044_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_8331_ _8331_/A _8331_/B vssd1 vssd1 vccd1 vccd1 _8331_/Y sky130_fd_sc_hd__nor2_1
X_5543_ _5578_/B _5542_/C _5542_/A vssd1 vssd1 vccd1 vccd1 _5554_/B sky130_fd_sc_hd__a21oi_1
X_8262_ _8262_/A _8262_/B vssd1 vssd1 vccd1 vccd1 _8495_/A sky130_fd_sc_hd__xnor2_1
X_5474_ _6034_/A _5879_/A vssd1 vssd1 vccd1 vccd1 _5514_/A sky130_fd_sc_hd__nand2_1
X_7213_ _7282_/A _7282_/B vssd1 vssd1 vccd1 vccd1 _7213_/X sky130_fd_sc_hd__or2b_1
X_8193_ _8398_/A vssd1 vssd1 vccd1 vccd1 _8194_/A sky130_fd_sc_hd__inv_2
X_4425_ _4426_/A vssd1 vssd1 vccd1 vccd1 _4425_/Y sky130_fd_sc_hd__inv_2
X_7144_ _7144_/A _7144_/B vssd1 vssd1 vccd1 vccd1 _7145_/B sky130_fd_sc_hd__xnor2_1
X_4356_ _4358_/A vssd1 vssd1 vccd1 vccd1 _4356_/Y sky130_fd_sc_hd__inv_2
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7075_ _7074_/A _7074_/B _7095_/A _7074_/D vssd1 vssd1 vccd1 vccd1 _7075_/X sky130_fd_sc_hd__o22a_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6026_ _6171_/B _6026_/B vssd1 vssd1 vccd1 vccd1 _6027_/B sky130_fd_sc_hd__xnor2_1
XFILLER_39_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7977_ _8022_/A _7976_/B _7976_/C vssd1 vssd1 vccd1 vccd1 _7978_/C sky130_fd_sc_hd__a21o_1
XFILLER_81_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6928_ _6737_/A _6737_/B _6839_/A _6839_/B _7092_/A vssd1 vssd1 vccd1 vccd1 _6977_/S
+ sky130_fd_sc_hd__a221o_1
XFILLER_42_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6859_ _7258_/A vssd1 vssd1 vccd1 vccd1 _7202_/A sky130_fd_sc_hd__buf_2
XFILLER_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8529_ _8533_/A _7583_/X _4650_/A vssd1 vssd1 vccd1 vccd1 _8529_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_89_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5190_ _5190_/A _5190_/B _5190_/C _5190_/D vssd1 vssd1 vccd1 vccd1 _5190_/X sky130_fd_sc_hd__or4_1
X_7900_ _7948_/A _7948_/B _7948_/C vssd1 vssd1 vccd1 vccd1 _7929_/A sky130_fd_sc_hd__nand3_1
XFILLER_55_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8880_ _8880_/A _4399_/Y vssd1 vssd1 vccd1 vccd1 io_out[27] sky130_fd_sc_hd__ebufn_8
XFILLER_36_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7831_ _7816_/A _7816_/B _7833_/B _7830_/A vssd1 vssd1 vccd1 vccd1 _7832_/B sky130_fd_sc_hd__a31o_1
XFILLER_51_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7762_ _7762_/A vssd1 vssd1 vccd1 vccd1 _8229_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_63_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4974_ _4979_/A vssd1 vssd1 vccd1 vccd1 _5174_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_7693_ _7693_/A _7693_/B vssd1 vssd1 vccd1 vccd1 _7745_/A sky130_fd_sc_hd__nor2_2
X_6713_ _6713_/A _6713_/B vssd1 vssd1 vccd1 vccd1 _6806_/B sky130_fd_sc_hd__xnor2_4
XFILLER_51_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6644_ _6614_/X _6642_/X _6643_/X _6798_/A _7238_/A vssd1 vssd1 vccd1 vccd1 _6718_/S
+ sky130_fd_sc_hd__a311o_4
X_6575_ _6581_/A _6581_/B vssd1 vssd1 vccd1 vccd1 _7176_/A sky130_fd_sc_hd__xor2_1
X_8314_ _8238_/A _8341_/B _8237_/B _8239_/B _8239_/A vssd1 vssd1 vccd1 vccd1 _8377_/A
+ sky130_fd_sc_hd__a32oi_4
X_5526_ _6323_/A _5879_/A _5526_/C vssd1 vssd1 vccd1 vccd1 _5526_/X sky130_fd_sc_hd__and3_1
X_8245_ _8455_/A _8245_/B vssd1 vssd1 vccd1 vccd1 _8292_/A sky130_fd_sc_hd__xnor2_1
X_5457_ _8662_/Q _7689_/B vssd1 vssd1 vccd1 vccd1 _5460_/A sky130_fd_sc_hd__nor2_2
X_4408_ _4408_/A vssd1 vssd1 vccd1 vccd1 _4408_/Y sky130_fd_sc_hd__inv_2
X_8176_ _8256_/B _8176_/B vssd1 vssd1 vccd1 vccd1 _8178_/B sky130_fd_sc_hd__xnor2_1
XFILLER_59_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5388_ _6364_/B vssd1 vssd1 vccd1 vccd1 _6371_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_7127_ _7425_/A _7030_/B _7032_/B _7035_/A vssd1 vssd1 vccd1 vccd1 _7128_/B sky130_fd_sc_hd__a31oi_2
X_4339_ _4339_/A vssd1 vssd1 vccd1 vccd1 _4339_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7058_ _7058_/A _7058_/B _7058_/C vssd1 vssd1 vccd1 vccd1 _7074_/A sky130_fd_sc_hd__and3_1
XFILLER_101_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6009_ _6009_/A _6215_/A vssd1 vssd1 vccd1 vccd1 _6009_/Y sky130_fd_sc_hd__nor2_1
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4690_ _5149_/A vssd1 vssd1 vccd1 vccd1 _5259_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6360_ _6358_/X _6359_/Y _5449_/B vssd1 vssd1 vccd1 vccd1 _6360_/Y sky130_fd_sc_hd__a21oi_1
X_5311_ input2/X _7545_/B vssd1 vssd1 vccd1 vccd1 _5320_/A sky130_fd_sc_hd__and2_1
X_8030_ _8030_/A _8109_/A vssd1 vssd1 vccd1 vccd1 _8031_/B sky130_fd_sc_hd__xnor2_1
X_6291_ _6192_/A _6192_/B _6193_/B _6193_/A vssd1 vssd1 vccd1 vccd1 _6294_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_102_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5242_ _5248_/B _5240_/X _5241_/X _5103_/B vssd1 vssd1 vccd1 vccd1 _5243_/D sky130_fd_sc_hd__o22a_1
X_5173_ _5214_/D _5173_/B _5176_/C _5173_/D vssd1 vssd1 vccd1 vccd1 _5173_/X sky130_fd_sc_hd__or4_1
XFILLER_68_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput1 active vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_6
XFILLER_96_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8863_ _8863_/A _4379_/Y vssd1 vssd1 vccd1 vccd1 io_out[10] sky130_fd_sc_hd__ebufn_8
X_7814_ _7814_/A _7814_/B vssd1 vssd1 vccd1 vccd1 _7815_/B sky130_fd_sc_hd__nand2_1
XFILLER_64_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7745_ _7745_/A _7745_/B vssd1 vssd1 vccd1 vccd1 _7864_/A sky130_fd_sc_hd__xor2_1
X_4957_ _5172_/A vssd1 vssd1 vccd1 vccd1 _5166_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7676_ _7676_/A _8713_/Q vssd1 vssd1 vccd1 vccd1 _7676_/X sky130_fd_sc_hd__or2b_1
X_4888_ _5135_/A vssd1 vssd1 vccd1 vccd1 _5143_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6627_ _6660_/A _6652_/B _6652_/C _6626_/Y vssd1 vssd1 vccd1 vccd1 _6657_/C sky130_fd_sc_hd__a31o_1
X_6558_ _6560_/B _8701_/Q vssd1 vssd1 vccd1 vccd1 _6710_/A sky130_fd_sc_hd__or2b_1
XFILLER_20_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6489_ _8704_/Q vssd1 vssd1 vccd1 vccd1 _7537_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_3_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5509_ _5482_/A _5508_/X _5506_/Y vssd1 vssd1 vccd1 vccd1 _5724_/C sky130_fd_sc_hd__a21o_1
X_8228_ _7885_/A _8326_/B _8406_/A _8406_/B vssd1 vssd1 vccd1 vccd1 _8334_/B sky130_fd_sc_hd__o22a_1
XFILLER_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8159_ _8254_/A _8159_/B vssd1 vssd1 vccd1 vccd1 _8161_/B sky130_fd_sc_hd__nor2_1
XFILLER_87_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5860_ _5862_/A _5862_/B vssd1 vssd1 vccd1 vccd1 _6074_/A sky130_fd_sc_hd__and2_1
XFILLER_34_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4811_ _4831_/A _4831_/B _4897_/B vssd1 vssd1 vccd1 vccd1 _4839_/B sky130_fd_sc_hd__or3_2
XFILLER_33_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5791_ _5895_/A vssd1 vssd1 vccd1 vccd1 _5997_/A sky130_fd_sc_hd__buf_2
X_7530_ _7526_/B _7527_/A _7526_/A vssd1 vssd1 vccd1 vccd1 _7532_/B sky130_fd_sc_hd__a21boi_1
X_4742_ _6406_/A vssd1 vssd1 vccd1 vccd1 _5296_/A sky130_fd_sc_hd__clkbuf_2
X_7461_ _7480_/A _7480_/B _7480_/C _7485_/B _7460_/X vssd1 vssd1 vccd1 vccd1 _7490_/B
+ sky130_fd_sc_hd__a41o_1
X_4673_ _4673_/A vssd1 vssd1 vccd1 vccd1 _4681_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6412_ _8666_/Q _8665_/Q _8667_/Q vssd1 vssd1 vccd1 vccd1 _6413_/B sky130_fd_sc_hd__a21o_1
X_7392_ _7305_/A _7320_/A _7306_/B _7220_/A vssd1 vssd1 vccd1 vccd1 _7396_/A sky130_fd_sc_hd__o2bb2ai_1
X_6343_ _5412_/A _5413_/A _6343_/S vssd1 vssd1 vccd1 vccd1 _6344_/A sky130_fd_sc_hd__mux2_1
X_6274_ _6274_/A _6274_/B vssd1 vssd1 vccd1 vccd1 _6297_/A sky130_fd_sc_hd__xnor2_2
X_8013_ _8013_/A _8017_/A _8013_/C vssd1 vssd1 vccd1 vccd1 _8015_/B sky130_fd_sc_hd__or3_1
X_5225_ _5223_/X _5224_/X _5060_/A vssd1 vssd1 vccd1 vccd1 _5261_/B sky130_fd_sc_hd__a21oi_1
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5156_ _5071_/A _4839_/B _4885_/X vssd1 vssd1 vccd1 vccd1 _5156_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_29_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5087_ _5087_/A _5243_/C vssd1 vssd1 vccd1 vccd1 _5087_/X sky130_fd_sc_hd__or2_1
XFILLER_84_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8915_ _8915_/A _4440_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[24] sky130_fd_sc_hd__ebufn_8
XFILLER_44_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8846_ _8846_/A _4358_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[25] sky130_fd_sc_hd__ebufn_8
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5989_ _6269_/A _6201_/B vssd1 vssd1 vccd1 vccd1 _5990_/B sky130_fd_sc_hd__xnor2_1
XFILLER_40_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7728_ _7853_/B _7777_/C _7727_/X vssd1 vssd1 vccd1 vccd1 _7729_/B sky130_fd_sc_hd__o21a_1
X_7659_ _7657_/X _7679_/A vssd1 vssd1 vccd1 vccd1 _7660_/B sky130_fd_sc_hd__and2b_1
XFILLER_4_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5010_ _5011_/A _5010_/B vssd1 vssd1 vccd1 vccd1 _5118_/B sky130_fd_sc_hd__nor2_2
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6961_ _6961_/A _6961_/B vssd1 vssd1 vccd1 vccd1 _6962_/B sky130_fd_sc_hd__xnor2_1
X_8700_ input3/X _8700_/D vssd1 vssd1 vccd1 vccd1 _8700_/Q sky130_fd_sc_hd__dfxtp_2
X_6892_ _6892_/A _6991_/A vssd1 vssd1 vccd1 vccd1 _6992_/A sky130_fd_sc_hd__xor2_1
XFILLER_81_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5912_ _6231_/A _5912_/B _5912_/C vssd1 vssd1 vccd1 vccd1 _5913_/B sky130_fd_sc_hd__and3_1
XFILLER_61_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8631_ input3/X _8631_/D vssd1 vssd1 vccd1 vccd1 _8631_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5843_ _5935_/B _5843_/B vssd1 vssd1 vccd1 vccd1 _5844_/B sky130_fd_sc_hd__nor2_1
X_8780__58 vssd1 vssd1 vccd1 vccd1 _8780__58/HI _8889_/A sky130_fd_sc_hd__conb_1
X_8562_ _8562_/A _8566_/B vssd1 vssd1 vccd1 vccd1 _8563_/B sky130_fd_sc_hd__nand2_1
XFILLER_34_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7513_ _8686_/Q _7514_/A vssd1 vssd1 vccd1 vccd1 _7515_/A sky130_fd_sc_hd__or2b_1
X_5774_ _6042_/B vssd1 vssd1 vccd1 vccd1 _5826_/B sky130_fd_sc_hd__inv_2
XFILLER_21_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8493_ _8493_/A _8493_/B vssd1 vssd1 vccd1 vccd1 _8493_/X sky130_fd_sc_hd__xor2_1
X_4725_ _4723_/A _5265_/A _4717_/A _4724_/X vssd1 vssd1 vccd1 vccd1 _8601_/D sky130_fd_sc_hd__o211a_1
X_7444_ _6589_/X _6596_/B _6590_/A vssd1 vssd1 vccd1 vccd1 _7495_/B sky130_fd_sc_hd__a21oi_1
X_4656_ _5245_/A vssd1 vssd1 vccd1 vccd1 _4657_/A sky130_fd_sc_hd__clkbuf_2
X_7375_ _7375_/A _7375_/B vssd1 vssd1 vccd1 vccd1 _7397_/A sky130_fd_sc_hd__xnor2_1
X_4587_ _4587_/A _4646_/A _4587_/C vssd1 vssd1 vccd1 vccd1 _4588_/A sky130_fd_sc_hd__and3_1
X_6326_ _6326_/A _6326_/B _6326_/C vssd1 vssd1 vccd1 vccd1 _6326_/X sky130_fd_sc_hd__or3_1
XFILLER_1_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6257_ _6257_/A _6257_/B vssd1 vssd1 vccd1 vccd1 _6260_/A sky130_fd_sc_hd__xnor2_1
XFILLER_57_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6188_ _6188_/A _6279_/B vssd1 vssd1 vccd1 vccd1 _6189_/B sky130_fd_sc_hd__xnor2_1
XFILLER_29_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5208_ _5190_/C _5207_/Y _4694_/A vssd1 vssd1 vccd1 vccd1 _5208_/X sky130_fd_sc_hd__o21a_1
XFILLER_69_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5139_ _5139_/A _5138_/Y vssd1 vssd1 vccd1 vccd1 _5139_/X sky130_fd_sc_hd__or2b_1
XFILLER_84_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8829_ _8829_/A _4337_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[8] sky130_fd_sc_hd__ebufn_8
XFILLER_40_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4510_ _7676_/A vssd1 vssd1 vccd1 vccd1 _5617_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5490_ _5881_/B _5533_/B vssd1 vssd1 vccd1 vccd1 _6034_/B sky130_fd_sc_hd__nand2_2
X_4441_ _4444_/A vssd1 vssd1 vccd1 vccd1 _4441_/Y sky130_fd_sc_hd__inv_2
X_7160_ _7219_/A _7160_/B vssd1 vssd1 vccd1 vccd1 _7161_/B sky130_fd_sc_hd__and2_1
X_4372_ _4396_/A vssd1 vssd1 vccd1 vccd1 _4377_/A sky130_fd_sc_hd__buf_6
X_6111_ _6044_/B _6125_/A _6111_/S vssd1 vssd1 vccd1 vccd1 _6113_/B sky130_fd_sc_hd__mux2_1
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7091_ _7087_/A _7087_/B _7090_/X vssd1 vssd1 vccd1 vccd1 _7158_/A sky130_fd_sc_hd__o21ai_2
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6042_ _6042_/A _6042_/B vssd1 vssd1 vccd1 vccd1 _6043_/A sky130_fd_sc_hd__nor2_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7993_ _8066_/A _7993_/B vssd1 vssd1 vccd1 vccd1 _8068_/B sky130_fd_sc_hd__and2b_1
X_6944_ _7060_/B _7135_/A vssd1 vssd1 vccd1 vccd1 _6944_/Y sky130_fd_sc_hd__nand2_1
XFILLER_54_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6875_ _6876_/B _6875_/B vssd1 vssd1 vccd1 vccd1 _7205_/B sky130_fd_sc_hd__xnor2_2
XFILLER_62_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8614_ input3/X _8614_/D vssd1 vssd1 vccd1 vccd1 _8614_/Q sky130_fd_sc_hd__dfxtp_1
X_5826_ _5826_/A _5826_/B vssd1 vssd1 vccd1 vccd1 _5870_/B sky130_fd_sc_hd__and2_1
XFILLER_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8545_ _8706_/Q vssd1 vssd1 vccd1 vccd1 _8561_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_5757_ _5850_/A _5756_/X vssd1 vssd1 vccd1 vccd1 _5824_/A sky130_fd_sc_hd__or2b_1
X_8476_ _8476_/A vssd1 vssd1 vccd1 vccd1 _8476_/Y sky130_fd_sc_hd__inv_2
X_4708_ _4705_/A _4697_/Y _4707_/X _4677_/X vssd1 vssd1 vccd1 vccd1 _8597_/D sky130_fd_sc_hd__o211a_1
X_7427_ _7428_/A _7428_/B vssd1 vssd1 vccd1 vccd1 _7434_/B sky130_fd_sc_hd__xnor2_1
X_5688_ _5688_/A _5688_/B vssd1 vssd1 vccd1 vccd1 _5710_/B sky130_fd_sc_hd__nand2_1
X_4639_ _4641_/B _4639_/B _4639_/C vssd1 vssd1 vccd1 vccd1 _4640_/A sky130_fd_sc_hd__and3b_1
X_7358_ _6765_/B _7320_/A _7220_/B _7306_/A vssd1 vssd1 vccd1 vccd1 _7368_/A sky130_fd_sc_hd__a22o_1
X_7289_ _7301_/A _7289_/B vssd1 vssd1 vccd1 vccd1 _7377_/A sky130_fd_sc_hd__xnor2_1
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6309_ _6309_/A _6309_/B vssd1 vssd1 vccd1 vccd1 _6326_/B sky130_fd_sc_hd__nor2_1
XFILLER_103_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4990_ _4990_/A _4990_/B vssd1 vssd1 vccd1 vccd1 _4990_/Y sky130_fd_sc_hd__nand2_1
XFILLER_44_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6660_ _6660_/A _6660_/B vssd1 vssd1 vccd1 vccd1 _6687_/A sky130_fd_sc_hd__nand2_1
X_8750__28 vssd1 vssd1 vccd1 vccd1 _8750__28/HI _8845_/A sky130_fd_sc_hd__conb_1
X_6591_ _6591_/A _6591_/B vssd1 vssd1 vccd1 vccd1 _7296_/A sky130_fd_sc_hd__nand2_2
X_5611_ _5657_/A _5657_/B vssd1 vssd1 vccd1 vccd1 _5671_/A sky130_fd_sc_hd__xnor2_1
X_8330_ _8334_/A vssd1 vssd1 vccd1 vccd1 _8407_/S sky130_fd_sc_hd__dlymetal6s2s_1
X_5542_ _5542_/A _5578_/B _5542_/C vssd1 vssd1 vccd1 vccd1 _5554_/A sky130_fd_sc_hd__and3_1
XFILLER_8_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8261_ _8428_/A _8428_/B vssd1 vssd1 vccd1 vccd1 _8262_/B sky130_fd_sc_hd__xor2_1
X_5473_ _5794_/A vssd1 vssd1 vccd1 vccd1 _5879_/A sky130_fd_sc_hd__clkbuf_2
X_7212_ _7212_/A _7212_/B vssd1 vssd1 vccd1 vccd1 _7282_/B sky130_fd_sc_hd__xnor2_1
X_4424_ _4426_/A vssd1 vssd1 vccd1 vccd1 _4424_/Y sky130_fd_sc_hd__inv_2
X_8192_ _8163_/A _8163_/B _8191_/Y vssd1 vssd1 vccd1 vccd1 _8272_/A sky130_fd_sc_hd__a21oi_1
X_7143_ _7018_/A _7018_/B _7142_/X vssd1 vssd1 vccd1 vccd1 _7144_/B sky130_fd_sc_hd__a21oi_1
X_4355_ _4358_/A vssd1 vssd1 vccd1 vccd1 _4355_/Y sky130_fd_sc_hd__inv_2
X_7074_ _7074_/A _7074_/B _7095_/A _7074_/D vssd1 vssd1 vccd1 vccd1 _7095_/B sky130_fd_sc_hd__nor4_2
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6025_ _6025_/A _6025_/B vssd1 vssd1 vccd1 vccd1 _6026_/B sky130_fd_sc_hd__xnor2_1
XFILLER_39_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7976_ _8022_/A _7976_/B _7976_/C vssd1 vssd1 vccd1 vccd1 _8022_/B sky130_fd_sc_hd__nand3_1
XFILLER_42_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6927_ _7160_/B _7031_/S vssd1 vssd1 vccd1 vccd1 _6931_/A sky130_fd_sc_hd__nor2_1
X_6858_ _7088_/B _6858_/B vssd1 vssd1 vccd1 vccd1 _7258_/A sky130_fd_sc_hd__and2_1
X_5809_ _5809_/A _5809_/B vssd1 vssd1 vccd1 vccd1 _5879_/C sky130_fd_sc_hd__xor2_1
X_6789_ _6789_/A _6722_/B vssd1 vssd1 vccd1 vccd1 _6823_/A sky130_fd_sc_hd__or2b_1
X_8528_ _4581_/A _8718_/Q _8514_/X _8527_/X vssd1 vssd1 vccd1 vccd1 _8718_/D sky130_fd_sc_hd__o22a_1
XFILLER_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8459_ _8326_/A _8406_/Y _7964_/X vssd1 vssd1 vccd1 vccd1 _8460_/B sky130_fd_sc_hd__o21ba_1
XFILLER_2_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7830_ _7830_/A _7830_/B vssd1 vssd1 vccd1 vccd1 _7833_/B sky130_fd_sc_hd__nor2_1
XFILLER_24_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7761_ _7764_/A _8111_/B _8111_/C vssd1 vssd1 vccd1 vccd1 _7762_/A sky130_fd_sc_hd__and3_1
X_4973_ _4990_/B _5017_/B vssd1 vssd1 vccd1 vccd1 _5004_/C sky130_fd_sc_hd__nand2_1
X_7692_ _8597_/Q _8539_/A vssd1 vssd1 vccd1 vccd1 _7693_/B sky130_fd_sc_hd__and2b_1
X_6712_ _6712_/A _6712_/B vssd1 vssd1 vccd1 vccd1 _6713_/B sky130_fd_sc_hd__nand2_2
X_6643_ _6657_/C vssd1 vssd1 vccd1 vccd1 _6643_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_32_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6574_ _8690_/Q _7634_/A vssd1 vssd1 vccd1 vccd1 _6581_/B sky130_fd_sc_hd__xnor2_2
X_8313_ _8313_/A _8313_/B vssd1 vssd1 vccd1 vccd1 _8376_/A sky130_fd_sc_hd__xnor2_1
X_5525_ _6034_/A vssd1 vssd1 vccd1 vccd1 _6323_/A sky130_fd_sc_hd__clkbuf_2
X_8244_ _8437_/A _8276_/B vssd1 vssd1 vccd1 vccd1 _8245_/B sky130_fd_sc_hd__xor2_1
X_5456_ _5881_/A vssd1 vssd1 vccd1 vccd1 _6034_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4407_ _4408_/A vssd1 vssd1 vccd1 vccd1 _4407_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_59_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8175_ _8079_/A _8079_/C _8079_/B vssd1 vssd1 vccd1 vccd1 _8176_/B sky130_fd_sc_hd__a21boi_1
X_5387_ _8664_/Q vssd1 vssd1 vccd1 vccd1 _5549_/A sky130_fd_sc_hd__inv_2
XFILLER_101_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7126_ _7012_/A _7012_/B _7011_/A vssd1 vssd1 vccd1 vccd1 _7128_/A sky130_fd_sc_hd__o21ai_1
X_4338_ _4339_/A vssd1 vssd1 vccd1 vccd1 _4338_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7057_ _7057_/A _7057_/B vssd1 vssd1 vccd1 vccd1 _7058_/C sky130_fd_sc_hd__nand2_1
XFILLER_86_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6008_ _6008_/A _6008_/B vssd1 vssd1 vccd1 vccd1 _6012_/B sky130_fd_sc_hd__xnor2_1
XFILLER_67_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7959_ _7958_/B _8025_/A _8117_/S vssd1 vssd1 vccd1 vccd1 _7960_/C sky130_fd_sc_hd__a21bo_1
XFILLER_42_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6290_ _6290_/A _6290_/B vssd1 vssd1 vccd1 vccd1 _6295_/A sky130_fd_sc_hd__xnor2_1
X_5310_ _8643_/Q _8642_/Q _5309_/X _8644_/Q vssd1 vssd1 vccd1 vccd1 _7545_/B sky130_fd_sc_hd__a31oi_4
X_5241_ _5241_/A _5241_/B _5241_/C vssd1 vssd1 vccd1 vccd1 _5241_/X sky130_fd_sc_hd__or3_1
XFILLER_96_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5172_ _5172_/A _5172_/B _5172_/C vssd1 vssd1 vccd1 vccd1 _5173_/D sky130_fd_sc_hd__or3_1
XFILLER_68_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput2 io_in[10] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__clkbuf_4
X_8862_ _8862_/A _4377_/Y vssd1 vssd1 vccd1 vccd1 io_out[9] sky130_fd_sc_hd__ebufn_8
XFILLER_64_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7813_ _7942_/B _7813_/B vssd1 vssd1 vccd1 vccd1 _7944_/A sky130_fd_sc_hd__nand2_1
XFILLER_64_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7744_ _8118_/A _7857_/C vssd1 vssd1 vccd1 vccd1 _7759_/A sky130_fd_sc_hd__xnor2_1
X_4956_ _5240_/B _4979_/A vssd1 vssd1 vccd1 vccd1 _5172_/A sky130_fd_sc_hd__or2_1
X_7675_ _7616_/A _7676_/A vssd1 vssd1 vccd1 vccd1 _7677_/A sky130_fd_sc_hd__and2b_1
XFILLER_20_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4887_ _4661_/A _4916_/B _5009_/B _4881_/X _4886_/X vssd1 vssd1 vccd1 vccd1 _4887_/X
+ sky130_fd_sc_hd__a2111o_1
X_6626_ _6626_/A _6664_/B vssd1 vssd1 vccd1 vccd1 _6626_/Y sky130_fd_sc_hd__nand2_1
X_6557_ _6592_/A _6584_/B _6556_/X vssd1 vssd1 vccd1 vccd1 _6562_/A sky130_fd_sc_hd__a21o_1
X_5508_ _5486_/A _5486_/B _5502_/Y vssd1 vssd1 vccd1 vccd1 _5508_/X sky130_fd_sc_hd__a21o_1
X_6488_ _8705_/Q _6505_/A _6488_/C vssd1 vssd1 vccd1 vccd1 _6488_/X sky130_fd_sc_hd__or3_1
X_8227_ _8120_/A _8225_/Y _8410_/A vssd1 vssd1 vccd1 vccd1 _8324_/A sky130_fd_sc_hd__o21a_1
X_5439_ _5413_/A _5436_/X _5442_/B _5412_/X _5447_/A vssd1 vssd1 vccd1 vccd1 _8651_/D
+ sky130_fd_sc_hd__a32o_1
X_8158_ _8158_/A _8158_/B vssd1 vssd1 vccd1 vccd1 _8159_/B sky130_fd_sc_hd__nor2_1
XFILLER_59_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7109_ _7236_/A _7197_/B vssd1 vssd1 vccd1 vccd1 _7110_/B sky130_fd_sc_hd__nand2_1
X_8089_ _8099_/B _8089_/B vssd1 vssd1 vccd1 vccd1 _8090_/B sky130_fd_sc_hd__xnor2_1
XFILLER_74_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8786__64 vssd1 vssd1 vccd1 vccd1 _8786__64/HI _8895_/A sky130_fd_sc_hd__conb_1
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4810_ _4810_/A _4810_/B vssd1 vssd1 vccd1 vccd1 _4897_/B sky130_fd_sc_hd__or2_2
XFILLER_61_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5790_ _5738_/A _5738_/B _5789_/Y vssd1 vssd1 vccd1 vccd1 _5815_/A sky130_fd_sc_hd__o21a_1
X_4741_ _4802_/B _4842_/C vssd1 vssd1 vccd1 vccd1 _4824_/C sky130_fd_sc_hd__nand2_1
X_7460_ _7459_/A _7367_/A _7459_/B vssd1 vssd1 vccd1 vccd1 _7460_/X sky130_fd_sc_hd__o21ba_1
X_4672_ _5243_/A _5105_/A vssd1 vssd1 vccd1 vccd1 _4673_/A sky130_fd_sc_hd__nor2_1
X_6411_ _8667_/Q _8666_/Q _8665_/Q vssd1 vssd1 vccd1 vccd1 _6416_/B sky130_fd_sc_hd__and3_1
X_7391_ _7393_/A _7393_/B vssd1 vssd1 vccd1 vccd1 _7395_/B sky130_fd_sc_hd__nor2_1
X_6342_ _6329_/X _6341_/X _6334_/X _8657_/Q vssd1 vssd1 vccd1 vccd1 _8657_/D sky130_fd_sc_hd__o2bb2a_1
XFILLER_88_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6273_ _6273_/A _6273_/B vssd1 vssd1 vccd1 vccd1 _6274_/B sky130_fd_sc_hd__xnor2_1
XFILLER_88_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8012_ _8019_/B _8010_/X _7938_/A _7940_/A vssd1 vssd1 vccd1 vccd1 _8013_/C sky130_fd_sc_hd__a211oi_1
X_5224_ _5259_/A _5259_/B _5224_/C _5224_/D vssd1 vssd1 vccd1 vccd1 _5224_/X sky130_fd_sc_hd__or4_1
XFILLER_96_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5155_ _5253_/B _5159_/C _5154_/X vssd1 vssd1 vccd1 vccd1 _5155_/X sky130_fd_sc_hd__or3b_1
X_5086_ _5086_/A vssd1 vssd1 vccd1 vccd1 _5243_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_84_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8914_ _8914_/A _4438_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[23] sky130_fd_sc_hd__ebufn_8
XFILLER_25_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8845_ _8845_/A _4357_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[24] sky130_fd_sc_hd__ebufn_8
XFILLER_71_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5988_ _5988_/A _5988_/B vssd1 vssd1 vccd1 vccd1 _6201_/B sky130_fd_sc_hd__xnor2_2
X_7727_ _8134_/A _8395_/B vssd1 vssd1 vccd1 vccd1 _7727_/X sky130_fd_sc_hd__or2_1
X_4939_ _4939_/A vssd1 vssd1 vccd1 vccd1 _5176_/C sky130_fd_sc_hd__clkbuf_2
X_7658_ _7658_/A _7658_/B vssd1 vssd1 vccd1 vccd1 _7679_/A sky130_fd_sc_hd__or2_1
XFILLER_20_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6609_ _6836_/A _6837_/A _6837_/B _6608_/X vssd1 vssd1 vccd1 vccd1 _6737_/B sky130_fd_sc_hd__a31o_2
X_7589_ _8708_/Q _7589_/B vssd1 vssd1 vccd1 vccd1 _7589_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6960_ _7004_/A _6960_/B vssd1 vssd1 vccd1 vccd1 _6961_/B sky130_fd_sc_hd__xnor2_1
XFILLER_81_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5911_ _6231_/A _5912_/B _5912_/C vssd1 vssd1 vccd1 vccd1 _5913_/A sky130_fd_sc_hd__a21oi_1
X_6891_ _7202_/A _6891_/B vssd1 vssd1 vccd1 vccd1 _6991_/A sky130_fd_sc_hd__xnor2_1
XFILLER_81_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8630_ input3/X _8630_/D vssd1 vssd1 vccd1 vccd1 _8630_/Q sky130_fd_sc_hd__dfxtp_1
X_5842_ _5842_/A _5842_/B vssd1 vssd1 vccd1 vccd1 _5843_/B sky130_fd_sc_hd__nor2_1
XFILLER_34_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8561_ _8561_/A _8561_/B vssd1 vssd1 vccd1 vccd1 _8566_/B sky130_fd_sc_hd__or2_1
X_5773_ _5954_/B _6284_/S _5974_/A vssd1 vssd1 vccd1 vccd1 _5777_/A sky130_fd_sc_hd__o21ai_1
X_7512_ _7512_/A vssd1 vssd1 vccd1 vccd1 _8699_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4724_ _4732_/A _4723_/X _4724_/S vssd1 vssd1 vccd1 vccd1 _4724_/X sky130_fd_sc_hd__mux2_1
X_8492_ _8492_/A _8492_/B _8492_/C vssd1 vssd1 vccd1 vccd1 _8492_/X sky130_fd_sc_hd__and3_1
X_7443_ _7443_/A _7443_/B vssd1 vssd1 vccd1 vccd1 _7495_/A sky130_fd_sc_hd__xnor2_1
X_4655_ _4989_/A vssd1 vssd1 vccd1 vccd1 _5245_/A sky130_fd_sc_hd__clkbuf_2
X_7374_ _7375_/A _7375_/B vssd1 vssd1 vccd1 vccd1 _7374_/X sky130_fd_sc_hd__or2b_1
X_4586_ _8572_/Q _8571_/Q vssd1 vssd1 vccd1 vccd1 _4587_/C sky130_fd_sc_hd__nand2_1
X_6325_ _6341_/A _6341_/B _6332_/A vssd1 vssd1 vccd1 vccd1 _6325_/X sky130_fd_sc_hd__or3_1
XFILLER_88_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6256_ _6227_/S _6226_/A _5587_/Y vssd1 vssd1 vccd1 vccd1 _6257_/B sky130_fd_sc_hd__a21o_1
X_6187_ _6187_/A _6187_/B vssd1 vssd1 vccd1 vccd1 _6279_/B sky130_fd_sc_hd__xor2_1
X_5207_ _4701_/A _5197_/X _5206_/X vssd1 vssd1 vccd1 vccd1 _5207_/Y sky130_fd_sc_hd__a21oi_1
X_5138_ _5214_/C _5138_/B _5239_/B _5199_/A vssd1 vssd1 vccd1 vccd1 _5138_/Y sky130_fd_sc_hd__nor4_1
XFILLER_96_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5069_ _5094_/B vssd1 vssd1 vccd1 vccd1 _5070_/D sky130_fd_sc_hd__clkbuf_2
X_8756__34 vssd1 vssd1 vccd1 vccd1 _8756__34/HI _8851_/A sky130_fd_sc_hd__conb_1
X_8828_ _8828_/A _4336_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[7] sky130_fd_sc_hd__ebufn_8
XFILLER_16_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4440_ _4444_/A vssd1 vssd1 vccd1 vccd1 _4440_/Y sky130_fd_sc_hd__inv_2
X_4371_ input1/X vssd1 vssd1 vccd1 vccd1 _4396_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_98_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6110_ _6123_/A _6110_/B vssd1 vssd1 vccd1 vccd1 _6111_/S sky130_fd_sc_hd__nand2_1
X_7090_ _7462_/B _7462_/A vssd1 vssd1 vccd1 vccd1 _7090_/X sky130_fd_sc_hd__or2b_1
XFILLER_98_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6041_ _6051_/B _6041_/B vssd1 vssd1 vccd1 vccd1 _6054_/A sky130_fd_sc_hd__xnor2_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7992_ _8006_/A _7992_/B _7996_/A vssd1 vssd1 vccd1 vccd1 _7993_/B sky130_fd_sc_hd__or3_1
XFILLER_66_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6943_ _6834_/A _6834_/B _6942_/X vssd1 vssd1 vccd1 vccd1 _6963_/A sky130_fd_sc_hd__o21ai_1
XFILLER_54_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6874_ _6883_/B _6876_/C _6876_/A vssd1 vssd1 vccd1 vccd1 _6875_/B sky130_fd_sc_hd__a21oi_1
X_5825_ _5962_/A _5961_/B vssd1 vssd1 vccd1 vccd1 _5983_/B sky130_fd_sc_hd__nor2b_2
X_8613_ input3/X _8613_/D vssd1 vssd1 vccd1 vccd1 _8613_/Q sky130_fd_sc_hd__dfxtp_1
X_8544_ _7581_/X _8542_/X _8543_/Y vssd1 vssd1 vccd1 vccd1 _8721_/D sky130_fd_sc_hd__o21a_1
X_5756_ _5959_/A _5755_/B _5755_/D _5755_/C vssd1 vssd1 vccd1 vccd1 _5756_/X sky130_fd_sc_hd__a31o_1
XFILLER_22_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8475_ _8475_/A _8475_/B vssd1 vssd1 vccd1 vccd1 _8479_/A sky130_fd_sc_hd__xnor2_1
X_5687_ _5688_/A _5688_/B vssd1 vssd1 vccd1 vccd1 _5768_/B sky130_fd_sc_hd__or2_1
X_4707_ _4707_/A _4707_/B vssd1 vssd1 vccd1 vccd1 _4707_/X sky130_fd_sc_hd__or2_1
X_7426_ _7424_/A _7424_/B _7431_/B _7431_/A vssd1 vssd1 vccd1 vccd1 _7428_/B sky130_fd_sc_hd__o22a_1
X_4638_ _8586_/Q _8587_/Q _4632_/B _8588_/Q vssd1 vssd1 vccd1 vccd1 _4639_/C sky130_fd_sc_hd__a31o_1
X_7357_ _7357_/A _7357_/B vssd1 vssd1 vccd1 vccd1 _7368_/B sky130_fd_sc_hd__xnor2_1
XFILLER_1_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4569_ input2/X vssd1 vssd1 vccd1 vccd1 _6406_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_103_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7288_ _7488_/A _7288_/B vssd1 vssd1 vccd1 vccd1 _7490_/A sky130_fd_sc_hd__nor2_1
XFILLER_89_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6308_ _6310_/A _6310_/B _6106_/A vssd1 vssd1 vccd1 vccd1 _6309_/B sky130_fd_sc_hd__a21o_1
X_6239_ _6239_/A _6275_/B vssd1 vssd1 vccd1 vccd1 _6240_/B sky130_fd_sc_hd__xnor2_2
XFILLER_76_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6590_ _6590_/A _6589_/X vssd1 vssd1 vccd1 vccd1 _6596_/A sky130_fd_sc_hd__or2b_1
X_5610_ _8648_/Q _7631_/B vssd1 vssd1 vccd1 vccd1 _5657_/B sky130_fd_sc_hd__xnor2_2
XFILLER_31_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5541_ _5881_/A _5540_/B _5540_/C _5578_/A vssd1 vssd1 vccd1 vccd1 _5542_/C sky130_fd_sc_hd__a22o_1
X_8260_ _8260_/A _8260_/B vssd1 vssd1 vccd1 vccd1 _8428_/B sky130_fd_sc_hd__xnor2_1
X_7211_ _7151_/A _7258_/B _7207_/B _7206_/B _7206_/A vssd1 vssd1 vccd1 vccd1 _7282_/A
+ sky130_fd_sc_hd__a32oi_4
X_5472_ _5486_/A _5486_/B vssd1 vssd1 vccd1 vccd1 _5794_/A sky130_fd_sc_hd__xor2_2
X_8191_ _8191_/A _8191_/B vssd1 vssd1 vccd1 vccd1 _8191_/Y sky130_fd_sc_hd__nor2_1
X_4423_ _4426_/A vssd1 vssd1 vccd1 vccd1 _4423_/Y sky130_fd_sc_hd__inv_2
X_7142_ _7017_/B _7142_/B vssd1 vssd1 vccd1 vccd1 _7142_/X sky130_fd_sc_hd__and2b_1
X_4354_ _4358_/A vssd1 vssd1 vccd1 vccd1 _4354_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7073_ _7072_/A _7072_/B _7072_/C vssd1 vssd1 vccd1 vccd1 _7074_/D sky130_fd_sc_hd__a21oi_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6024_ _6024_/A _6175_/B vssd1 vssd1 vccd1 vccd1 _6025_/B sky130_fd_sc_hd__xnor2_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7975_ _8044_/A _7975_/B vssd1 vssd1 vccd1 vccd1 _7976_/C sky130_fd_sc_hd__xnor2_1
XFILLER_27_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6926_ _6925_/A _6925_/B _6925_/C vssd1 vssd1 vccd1 vccd1 _6932_/B sky130_fd_sc_hd__a21o_1
XFILLER_54_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6857_ _7220_/A _7092_/C vssd1 vssd1 vccd1 vccd1 _6858_/B sky130_fd_sc_hd__nand2_1
X_6788_ _7190_/A _7190_/B _6735_/A vssd1 vssd1 vccd1 vccd1 _6854_/A sky130_fd_sc_hd__a21o_1
XFILLER_50_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5808_ _5898_/A _5895_/B vssd1 vssd1 vccd1 vccd1 _5809_/B sky130_fd_sc_hd__xnor2_1
X_8527_ _8527_/A _8527_/B _8527_/C vssd1 vssd1 vccd1 vccd1 _8527_/X sky130_fd_sc_hd__and3_1
X_5739_ _5739_/A _5739_/B vssd1 vssd1 vccd1 vccd1 _5744_/A sky130_fd_sc_hd__xor2_2
XFILLER_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8458_ _7766_/A _7766_/C _7871_/X vssd1 vssd1 vccd1 vccd1 _8460_/A sky130_fd_sc_hd__a21o_1
X_8389_ _8389_/A _8389_/B vssd1 vssd1 vccd1 vccd1 _8390_/B sky130_fd_sc_hd__nor2_1
X_7409_ _7409_/A _7409_/B _7409_/C vssd1 vssd1 vccd1 vccd1 _7413_/A sky130_fd_sc_hd__nand3_1
XFILLER_89_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8810__88 vssd1 vssd1 vccd1 vccd1 _8810__88/HI _8919_/A sky130_fd_sc_hd__conb_1
XFILLER_63_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7760_ _7760_/A _7853_/C vssd1 vssd1 vccd1 vccd1 _7772_/A sky130_fd_sc_hd__xnor2_1
X_4972_ _5119_/B _5072_/B vssd1 vssd1 vccd1 vccd1 _5017_/B sky130_fd_sc_hd__nor2_1
XFILLER_24_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7691_ _8721_/Q _8597_/Q vssd1 vssd1 vccd1 vccd1 _7693_/A sky130_fd_sc_hd__and2b_1
X_6711_ _6711_/A _6605_/B vssd1 vssd1 vccd1 vccd1 _6712_/B sky130_fd_sc_hd__or2b_1
X_6642_ _6657_/B vssd1 vssd1 vccd1 vccd1 _6642_/X sky130_fd_sc_hd__clkbuf_2
X_8312_ _8312_/A _8312_/B vssd1 vssd1 vccd1 vccd1 _8313_/B sky130_fd_sc_hd__xor2_1
X_6573_ _6591_/A _6580_/B _6572_/X vssd1 vssd1 vccd1 vccd1 _6581_/A sky130_fd_sc_hd__a21o_1
X_5524_ _6082_/B _5906_/A _5524_/C vssd1 vssd1 vccd1 vccd1 _6033_/B sky130_fd_sc_hd__and3_1
X_8243_ _8363_/A _8146_/B _8196_/X vssd1 vssd1 vccd1 vccd1 _8276_/B sky130_fd_sc_hd__o21a_1
X_5455_ _5584_/A _5534_/B vssd1 vssd1 vccd1 vccd1 _5881_/A sky130_fd_sc_hd__xor2_2
X_4406_ _4408_/A vssd1 vssd1 vccd1 vccd1 _4406_/Y sky130_fd_sc_hd__inv_2
X_8174_ _8172_/Y _8174_/B vssd1 vssd1 vccd1 vccd1 _8256_/B sky130_fd_sc_hd__and2b_1
XFILLER_99_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7125_ _7078_/B _7081_/A _7123_/Y _7124_/Y vssd1 vssd1 vccd1 vccd1 _7146_/A sky130_fd_sc_hd__o31a_2
X_5386_ _8664_/Q _5402_/C _5381_/X _5385_/X vssd1 vssd1 vccd1 vccd1 _5386_/X sky130_fd_sc_hd__o31a_1
XFILLER_101_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4337_ _4339_/A vssd1 vssd1 vccd1 vccd1 _4337_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7056_ _7052_/A _7101_/B _7055_/C vssd1 vssd1 vccd1 vccd1 _7058_/B sky130_fd_sc_hd__a21o_1
XFILLER_75_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6007_ _6007_/A _6007_/B vssd1 vssd1 vccd1 vccd1 _6008_/B sky130_fd_sc_hd__xor2_1
XFILLER_55_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7958_ _8117_/S _7958_/B _8025_/A vssd1 vssd1 vccd1 vccd1 _8025_/B sky130_fd_sc_hd__nand3b_1
XFILLER_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7889_ _7889_/A _7963_/A vssd1 vssd1 vccd1 vccd1 _7890_/B sky130_fd_sc_hd__nand2_1
X_6909_ _7135_/A _7057_/A _6909_/C vssd1 vssd1 vccd1 vccd1 _7057_/B sky130_fd_sc_hd__nand3_1
XFILLER_6_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5240_ _5240_/A _5240_/B _5240_/C _5237_/Y vssd1 vssd1 vccd1 vccd1 _5240_/X sky130_fd_sc_hd__or4b_1
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5171_ _4928_/Y _5135_/X _5253_/A vssd1 vssd1 vccd1 vccd1 _5171_/X sky130_fd_sc_hd__o21a_1
XFILLER_96_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput3 wb_clk_i vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_16
XFILLER_49_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8861_ _8861_/A _4376_/Y vssd1 vssd1 vccd1 vccd1 io_out[8] sky130_fd_sc_hd__ebufn_8
XFILLER_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7812_ _7812_/A _7812_/B vssd1 vssd1 vccd1 vccd1 _7813_/B sky130_fd_sc_hd__nand2_1
XFILLER_24_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7743_ _7758_/A _7743_/B vssd1 vssd1 vccd1 vccd1 _7857_/C sky130_fd_sc_hd__xnor2_1
X_4955_ _5011_/A _4955_/B vssd1 vssd1 vccd1 vccd1 _4979_/A sky130_fd_sc_hd__nor2_1
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7674_ _7788_/A vssd1 vssd1 vccd1 vccd1 _7904_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4886_ _5075_/B _4823_/B _5026_/C _4885_/X vssd1 vssd1 vccd1 vccd1 _4886_/X sky130_fd_sc_hd__a31o_1
XFILLER_32_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6625_ _8693_/Q _8610_/Q vssd1 vssd1 vccd1 vccd1 _6664_/B sky130_fd_sc_hd__or2b_1
X_6556_ _8700_/Q _6556_/B vssd1 vssd1 vccd1 vccd1 _6556_/X sky130_fd_sc_hd__and2b_1
X_5507_ _5507_/A _5507_/B _5506_/Y vssd1 vssd1 vccd1 vccd1 _5724_/B sky130_fd_sc_hd__or3b_2
X_8226_ _8226_/A vssd1 vssd1 vccd1 vccd1 _8410_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6487_ _7518_/B _7514_/A _6711_/A vssd1 vssd1 vccd1 vccd1 _6488_/C sky130_fd_sc_hd__o21a_1
X_5438_ _5448_/S vssd1 vssd1 vccd1 vccd1 _5442_/B sky130_fd_sc_hd__inv_2
X_8157_ _8158_/A _8158_/B vssd1 vssd1 vccd1 vccd1 _8254_/A sky130_fd_sc_hd__and2_1
X_5369_ _8641_/Q _5369_/B vssd1 vssd1 vccd1 vccd1 _5373_/B sky130_fd_sc_hd__and2_1
X_8088_ _8088_/A _8088_/B vssd1 vssd1 vccd1 vccd1 _8089_/B sky130_fd_sc_hd__xnor2_1
X_7108_ _6839_/A _6839_/B _7193_/A vssd1 vssd1 vccd1 vccd1 _7195_/A sky130_fd_sc_hd__a21o_1
X_7039_ _7039_/A _7039_/B vssd1 vssd1 vccd1 vccd1 _7039_/Y sky130_fd_sc_hd__nor2_1
XFILLER_74_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4740_ _4760_/A vssd1 vssd1 vccd1 vccd1 _5275_/B sky130_fd_sc_hd__clkbuf_2
X_4671_ _5183_/S vssd1 vssd1 vccd1 vccd1 _5105_/A sky130_fd_sc_hd__clkbuf_2
X_7390_ _7390_/A _7390_/B vssd1 vssd1 vccd1 vccd1 _7393_/B sky130_fd_sc_hd__xnor2_1
X_6410_ _6410_/A vssd1 vssd1 vccd1 vccd1 _8666_/D sky130_fd_sc_hd__clkbuf_1
X_6341_ _6341_/A _6341_/B _6340_/X vssd1 vssd1 vccd1 vccd1 _6341_/X sky130_fd_sc_hd__or3b_1
X_6272_ _6272_/A _6272_/B vssd1 vssd1 vccd1 vccd1 _6273_/B sky130_fd_sc_hd__xnor2_1
X_8011_ _7938_/A _7940_/A _8019_/B _8010_/X vssd1 vssd1 vccd1 vccd1 _8017_/A sky130_fd_sc_hd__o211a_1
X_5223_ _5251_/A _5223_/B vssd1 vssd1 vccd1 vccd1 _5223_/X sky130_fd_sc_hd__or2_1
X_5154_ _5214_/A _5152_/Y _5153_/Y _4886_/X _5057_/A vssd1 vssd1 vccd1 vccd1 _5154_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_96_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5085_ _5119_/A _5248_/A _5122_/B vssd1 vssd1 vccd1 vccd1 _5252_/B sky130_fd_sc_hd__or3_1
X_8913_ _8913_/A _4437_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[22] sky130_fd_sc_hd__ebufn_8
XFILLER_56_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8844_ _8844_/A _4356_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[23] sky130_fd_sc_hd__ebufn_8
XFILLER_71_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5987_ _6203_/A _5985_/A _6277_/B _6178_/A vssd1 vssd1 vccd1 vccd1 _5988_/B sky130_fd_sc_hd__o22a_1
X_7726_ _8116_/C _8116_/B vssd1 vssd1 vccd1 vccd1 _8395_/B sky130_fd_sc_hd__nand2_1
X_4938_ _4969_/C vssd1 vssd1 vccd1 vccd1 _5173_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_7657_ _7658_/A _8609_/Q vssd1 vssd1 vccd1 vccd1 _7657_/X sky130_fd_sc_hd__and2_1
X_4869_ _5219_/C _5030_/C vssd1 vssd1 vccd1 vccd1 _5023_/A sky130_fd_sc_hd__or2_1
X_6608_ _7537_/A _6608_/B vssd1 vssd1 vccd1 vccd1 _6608_/X sky130_fd_sc_hd__and2b_1
X_7588_ _7588_/A _7588_/B vssd1 vssd1 vccd1 vccd1 _7589_/B sky130_fd_sc_hd__nand2_1
X_6539_ _6539_/A _8687_/Q vssd1 vssd1 vccd1 vccd1 _6540_/D sky130_fd_sc_hd__or2_1
XFILLER_97_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8209_ _8209_/A _8462_/B vssd1 vssd1 vccd1 vccd1 _8381_/A sky130_fd_sc_hd__nand2_1
XFILLER_47_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5910_ _6017_/B _5910_/B vssd1 vssd1 vccd1 vccd1 _5912_/C sky130_fd_sc_hd__nand2_1
X_6890_ _6968_/B _6890_/B vssd1 vssd1 vccd1 vccd1 _6891_/B sky130_fd_sc_hd__xnor2_1
XFILLER_34_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5841_ _5842_/A _5842_/B vssd1 vssd1 vccd1 vccd1 _5935_/B sky130_fd_sc_hd__and2_1
XFILLER_34_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8560_ _8561_/A _8561_/B vssd1 vssd1 vccd1 vccd1 _8562_/A sky130_fd_sc_hd__nand2_1
X_5772_ _6063_/A _6063_/B vssd1 vssd1 vccd1 vccd1 _5781_/A sky130_fd_sc_hd__and2_1
X_8491_ _8492_/B _8492_/C _8492_/A vssd1 vssd1 vccd1 vccd1 _8491_/Y sky130_fd_sc_hd__a21oi_1
X_7511_ _6511_/A _6512_/A _7511_/S vssd1 vssd1 vccd1 vccd1 _7512_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4723_ _4723_/A _5265_/A vssd1 vssd1 vccd1 vccd1 _4723_/X sky130_fd_sc_hd__or2b_1
X_7442_ _7442_/A _7442_/B vssd1 vssd1 vccd1 vccd1 _7494_/A sky130_fd_sc_hd__xnor2_2
X_4654_ _5180_/A vssd1 vssd1 vccd1 vccd1 _4989_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7373_ _7373_/A _7373_/B vssd1 vssd1 vccd1 vccd1 _7375_/B sky130_fd_sc_hd__xor2_1
X_4585_ _4607_/A vssd1 vssd1 vccd1 vccd1 _4646_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6324_ _6327_/A _6322_/X _6323_/X vssd1 vssd1 vccd1 vccd1 _6332_/A sky130_fd_sc_hd__a21oi_1
X_6255_ _5482_/A _5508_/X _5546_/X vssd1 vssd1 vccd1 vccd1 _6257_/A sky130_fd_sc_hd__a21oi_2
X_5206_ _5199_/Y _5200_/X _5205_/Y _4995_/A vssd1 vssd1 vccd1 vccd1 _5206_/X sky130_fd_sc_hd__o211a_1
XFILLER_69_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6186_ _6186_/A _6281_/B vssd1 vssd1 vccd1 vccd1 _6187_/B sky130_fd_sc_hd__xnor2_1
X_5137_ _5151_/A _5137_/B _5137_/C vssd1 vssd1 vccd1 vccd1 _5137_/X sky130_fd_sc_hd__or3_1
X_5068_ _5068_/A _8592_/Q vssd1 vssd1 vccd1 vccd1 _5094_/B sky130_fd_sc_hd__nand2_1
XFILLER_84_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8827_ _8827_/A _4335_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[6] sky130_fd_sc_hd__ebufn_8
XFILLER_13_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8771__49 vssd1 vssd1 vccd1 vccd1 _8771__49/HI _8880_/A sky130_fd_sc_hd__conb_1
X_7709_ _7722_/A _7714_/B vssd1 vssd1 vccd1 vccd1 _7823_/A sky130_fd_sc_hd__nand2_1
X_8689_ input3/X _8689_/D vssd1 vssd1 vccd1 vccd1 _8689_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_79_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4370_ _4370_/A vssd1 vssd1 vccd1 vccd1 _4370_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6040_ _6040_/A _6040_/B vssd1 vssd1 vccd1 vccd1 _6057_/A sky130_fd_sc_hd__xnor2_1
XFILLER_100_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7991_ _8006_/A _7992_/B _7996_/A vssd1 vssd1 vccd1 vccd1 _8066_/A sky130_fd_sc_hd__o21a_1
XFILLER_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6942_ _6942_/A _6942_/B vssd1 vssd1 vccd1 vccd1 _6942_/X sky130_fd_sc_hd__or2_1
X_6873_ _7226_/B vssd1 vssd1 vccd1 vccd1 _6876_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_62_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5824_ _5824_/A _5824_/B vssd1 vssd1 vccd1 vccd1 _5842_/A sky130_fd_sc_hd__nor2_1
X_8612_ input3/X _8612_/D vssd1 vssd1 vccd1 vccd1 _8612_/Q sky130_fd_sc_hd__dfxtp_1
X_8543_ _8538_/A _7583_/X _4650_/A vssd1 vssd1 vccd1 vccd1 _8543_/Y sky130_fd_sc_hd__a21oi_1
X_5755_ _5959_/A _5755_/B _5755_/C _5755_/D vssd1 vssd1 vccd1 vccd1 _5850_/A sky130_fd_sc_hd__and4_1
X_8474_ _8390_/A _8390_/B _8389_/A vssd1 vssd1 vccd1 vccd1 _8475_/B sky130_fd_sc_hd__a21o_1
X_5686_ _6180_/A _5675_/B _5682_/A _5682_/B _5685_/Y vssd1 vssd1 vccd1 vccd1 _5688_/B
+ sky130_fd_sc_hd__o41a_1
XFILLER_30_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4706_ _5127_/A _5127_/B vssd1 vssd1 vccd1 vccd1 _4707_/B sky130_fd_sc_hd__nor2_1
X_7425_ _7425_/A _7425_/B vssd1 vssd1 vccd1 vccd1 _7431_/A sky130_fd_sc_hd__nand2_1
X_4637_ _8588_/Q _8587_/Q _4637_/C vssd1 vssd1 vccd1 vccd1 _4641_/B sky130_fd_sc_hd__and3_1
X_7356_ _7357_/A _7357_/B vssd1 vssd1 vccd1 vccd1 _7366_/B sky130_fd_sc_hd__nand2_1
X_4568_ _4568_/A vssd1 vssd1 vccd1 vccd1 _8873_/A sky130_fd_sc_hd__clkbuf_1
X_7287_ _7287_/A _7287_/B vssd1 vssd1 vccd1 vccd1 _7288_/B sky130_fd_sc_hd__and2_1
X_4499_ _8603_/Q vssd1 vssd1 vccd1 vccd1 _4810_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6307_ _6307_/A _6307_/B vssd1 vssd1 vccd1 vccd1 _6309_/A sky130_fd_sc_hd__xnor2_1
XFILLER_89_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6238_ _6238_/A _6238_/B vssd1 vssd1 vccd1 vccd1 _6275_/B sky130_fd_sc_hd__xor2_1
X_8816__94 vssd1 vssd1 vccd1 vccd1 _8816__94/HI _8925_/A sky130_fd_sc_hd__conb_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6169_ _6076_/Y _6310_/A _6310_/B _6168_/X vssd1 vssd1 vccd1 vccd1 _6306_/B sky130_fd_sc_hd__a31o_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5540_ _5881_/A _5540_/B _5540_/C _5578_/A vssd1 vssd1 vccd1 vccd1 _5578_/B sky130_fd_sc_hd__nand4_1
XFILLER_8_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5471_ _5475_/A _5475_/B _5477_/B _5470_/X _5468_/A vssd1 vssd1 vccd1 vccd1 _5486_/B
+ sky130_fd_sc_hd__a311o_4
X_7210_ _7212_/B _7212_/A vssd1 vssd1 vccd1 vccd1 _7210_/X sky130_fd_sc_hd__or2b_1
X_4422_ _4426_/A vssd1 vssd1 vccd1 vccd1 _4422_/Y sky130_fd_sc_hd__inv_2
X_8190_ _8181_/A _8181_/B _8189_/X vssd1 vssd1 vccd1 vccd1 _8269_/A sky130_fd_sc_hd__a21boi_1
X_4353_ _4365_/A vssd1 vssd1 vccd1 vccd1 _4358_/A sky130_fd_sc_hd__buf_2
X_7141_ _7141_/A _7141_/B vssd1 vssd1 vccd1 vccd1 _7144_/A sky130_fd_sc_hd__xnor2_1
X_7072_ _7072_/A _7072_/B _7072_/C vssd1 vssd1 vccd1 vccd1 _7095_/A sky130_fd_sc_hd__and3_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6023_ _6198_/A _6023_/B vssd1 vssd1 vccd1 vccd1 _6175_/B sky130_fd_sc_hd__xnor2_1
XFILLER_100_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7974_ _8043_/A _8043_/B vssd1 vssd1 vccd1 vccd1 _7975_/B sky130_fd_sc_hd__xor2_1
XFILLER_66_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6925_ _6925_/A _6925_/B _6925_/C vssd1 vssd1 vccd1 vccd1 _6932_/A sky130_fd_sc_hd__nand3_1
X_6856_ _7265_/B vssd1 vssd1 vccd1 vccd1 _7220_/A sky130_fd_sc_hd__buf_2
XFILLER_80_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6787_ _6787_/A _6787_/B vssd1 vssd1 vccd1 vccd1 _7190_/B sky130_fd_sc_hd__xor2_1
X_8741__19 vssd1 vssd1 vccd1 vccd1 _8741__19/HI _8836_/A sky130_fd_sc_hd__conb_1
XFILLER_10_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5807_ _5879_/A _5896_/A vssd1 vssd1 vccd1 vccd1 _5810_/A sky130_fd_sc_hd__nand2_1
X_8526_ _7845_/A _7847_/A _8526_/S vssd1 vssd1 vccd1 vccd1 _8527_/C sky130_fd_sc_hd__mux2_1
X_5738_ _5738_/A _5738_/B vssd1 vssd1 vccd1 vccd1 _5739_/B sky130_fd_sc_hd__xnor2_2
XFILLER_50_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8457_ _8403_/A _8403_/B _8401_/A vssd1 vssd1 vccd1 vccd1 _8465_/A sky130_fd_sc_hd__o21a_1
XFILLER_89_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5669_ _5826_/A vssd1 vssd1 vccd1 vccd1 _5754_/A sky130_fd_sc_hd__clkbuf_2
X_8388_ _8388_/A _8388_/B _8388_/C vssd1 vssd1 vccd1 vccd1 _8389_/B sky130_fd_sc_hd__and3_1
X_7408_ _7388_/A _7388_/C _7388_/B vssd1 vssd1 vccd1 vccd1 _7409_/C sky130_fd_sc_hd__o21ai_1
X_7339_ _7339_/A _7339_/B vssd1 vssd1 vccd1 vccd1 _7343_/A sky130_fd_sc_hd__nand2_1
XFILLER_104_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4971_ _5138_/B _5193_/B vssd1 vssd1 vccd1 vccd1 _5091_/D sky130_fd_sc_hd__or2_1
X_7690_ _7747_/A _7690_/B vssd1 vssd1 vccd1 vccd1 _7740_/A sky130_fd_sc_hd__nor2_4
X_6710_ _6710_/A _6710_/B vssd1 vssd1 vccd1 vccd1 _6713_/A sky130_fd_sc_hd__nand2_2
XFILLER_44_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6641_ _7418_/A _7020_/A vssd1 vssd1 vccd1 vccd1 _6641_/X sky130_fd_sc_hd__or2_1
X_8311_ _8385_/A _8379_/B vssd1 vssd1 vccd1 vccd1 _8312_/B sky130_fd_sc_hd__xnor2_1
X_6572_ _8689_/Q _8606_/Q vssd1 vssd1 vccd1 vccd1 _6572_/X sky130_fd_sc_hd__and2b_1
X_5523_ _6005_/A _6006_/A vssd1 vssd1 vccd1 vccd1 _5524_/C sky130_fd_sc_hd__nand2_1
X_8242_ _8272_/A _8272_/B vssd1 vssd1 vccd1 vccd1 _8258_/A sky130_fd_sc_hd__xor2_1
X_5454_ _8659_/Q _8596_/Q vssd1 vssd1 vccd1 vccd1 _5534_/B sky130_fd_sc_hd__xnor2_4
X_4405_ _4408_/A vssd1 vssd1 vccd1 vccd1 _4405_/Y sky130_fd_sc_hd__inv_2
X_8173_ _8172_/A _8172_/C _8172_/B vssd1 vssd1 vccd1 vccd1 _8174_/B sky130_fd_sc_hd__o21ai_1
X_5385_ _5462_/B _6346_/A _8658_/Q _5384_/Y vssd1 vssd1 vccd1 vccd1 _5385_/X sky130_fd_sc_hd__a31o_1
X_7124_ _7078_/B _7081_/A _7123_/Y vssd1 vssd1 vccd1 vccd1 _7124_/Y sky130_fd_sc_hd__o21ai_1
X_4336_ _4339_/A vssd1 vssd1 vccd1 vccd1 _4336_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7055_ _7115_/B _7101_/B _7055_/C vssd1 vssd1 vccd1 vccd1 _7058_/A sky130_fd_sc_hd__nand3_1
XFILLER_101_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6006_ _6006_/A _6224_/A vssd1 vssd1 vccd1 vccd1 _6007_/B sky130_fd_sc_hd__xnor2_1
XFILLER_27_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7957_ _7957_/A _8326_/A _7957_/C _7957_/D vssd1 vssd1 vccd1 vccd1 _8025_/A sky130_fd_sc_hd__or4_1
X_7888_ _7889_/A _7963_/A vssd1 vssd1 vccd1 vccd1 _8044_/A sky130_fd_sc_hd__or2_1
X_6908_ _6907_/B _6907_/C _7045_/A vssd1 vssd1 vccd1 vccd1 _6909_/C sky130_fd_sc_hd__a21bo_1
X_6839_ _6839_/A _6839_/B vssd1 vssd1 vccd1 vccd1 _6864_/A sky130_fd_sc_hd__and2_1
XFILLER_24_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8509_ _7664_/A _7816_/B _7887_/A _7853_/B _8508_/X vssd1 vssd1 vccd1 vccd1 _8520_/A
+ sky130_fd_sc_hd__a41o_1
XFILLER_2_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5170_ _5165_/X _5169_/X _5139_/A vssd1 vssd1 vccd1 vccd1 _5170_/X sky130_fd_sc_hd__a21o_1
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8860_ _8860_/A _4375_/Y vssd1 vssd1 vccd1 vccd1 io_out[7] sky130_fd_sc_hd__ebufn_8
XFILLER_91_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7811_ _7812_/A _7812_/B vssd1 vssd1 vccd1 vccd1 _7942_/B sky130_fd_sc_hd__or2_1
X_7742_ _7862_/A _7957_/A _8116_/B _7741_/Y vssd1 vssd1 vccd1 vccd1 _7743_/B sky130_fd_sc_hd__o211a_1
X_4954_ _4728_/B _4942_/X _4951_/X _4953_/X vssd1 vssd1 vccd1 vccd1 _4954_/X sky130_fd_sc_hd__o31a_1
XFILLER_51_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7673_ _7673_/A _7673_/B vssd1 vssd1 vccd1 vccd1 _7788_/A sky130_fd_sc_hd__or2_1
X_4885_ _5194_/A vssd1 vssd1 vccd1 vccd1 _4885_/X sky130_fd_sc_hd__clkbuf_2
X_6624_ _6626_/A _6624_/B vssd1 vssd1 vccd1 vccd1 _6652_/C sky130_fd_sc_hd__and2_1
X_6555_ _8700_/Q _6556_/B vssd1 vssd1 vccd1 vccd1 _6584_/B sky130_fd_sc_hd__xnor2_4
XFILLER_3_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5506_ _5506_/A _5506_/B vssd1 vssd1 vccd1 vccd1 _5506_/Y sky130_fd_sc_hd__nor2_1
X_8225_ _8225_/A _8319_/A vssd1 vssd1 vccd1 vccd1 _8225_/Y sky130_fd_sc_hd__nor2_1
X_6486_ _7518_/B _7514_/A _8699_/Q _7526_/A vssd1 vssd1 vccd1 vccd1 _6486_/X sky130_fd_sc_hd__a31o_1
X_5437_ _5442_/A _5437_/B _5437_/C vssd1 vssd1 vccd1 vccd1 _5448_/S sky130_fd_sc_hd__and3_1
XFILLER_99_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8156_ _8202_/A _8156_/B vssd1 vssd1 vccd1 vccd1 _8158_/B sky130_fd_sc_hd__and2_1
XFILLER_86_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5368_ _5369_/B _5368_/B vssd1 vssd1 vccd1 vccd1 _8640_/D sky130_fd_sc_hd__nor2_1
XFILLER_101_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8087_ _8185_/A _8087_/B vssd1 vssd1 vccd1 vccd1 _8088_/B sky130_fd_sc_hd__and2_1
X_7107_ _7107_/A _7137_/B vssd1 vssd1 vccd1 vccd1 _7107_/Y sky130_fd_sc_hd__nand2_1
X_5299_ _8697_/Q _5285_/A _5298_/X _5296_/X vssd1 vssd1 vccd1 vccd1 _8622_/D sky130_fd_sc_hd__o211a_1
XFILLER_101_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7038_ _7039_/A _7039_/B vssd1 vssd1 vccd1 vccd1 _7038_/Y sky130_fd_sc_hd__nand2_1
XFILLER_19_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8777__55 vssd1 vssd1 vccd1 vccd1 _8777__55/HI _8886_/A sky130_fd_sc_hd__conb_1
XFILLER_73_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4670_ _5235_/A vssd1 vssd1 vccd1 vccd1 _5183_/S sky130_fd_sc_hd__clkbuf_2
X_6340_ _6300_/A _6301_/X _6340_/S vssd1 vssd1 vccd1 vccd1 _6340_/X sky130_fd_sc_hd__mux2_1
X_6271_ _6271_/A _6271_/B vssd1 vssd1 vccd1 vccd1 _6272_/B sky130_fd_sc_hd__xnor2_1
X_8010_ _8019_/A _8009_/B _8009_/C vssd1 vssd1 vccd1 vccd1 _8010_/X sky130_fd_sc_hd__a21o_1
X_5222_ _4728_/B _5190_/C _5217_/X _5221_/X _5259_/A vssd1 vssd1 vccd1 vccd1 _5223_/B
+ sky130_fd_sc_hd__o32a_1
XFILLER_102_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5153_ _5153_/A _5153_/B vssd1 vssd1 vccd1 vccd1 _5153_/Y sky130_fd_sc_hd__nor2_1
XFILLER_69_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5084_ _5075_/B _5253_/C _5135_/C _5083_/X vssd1 vssd1 vccd1 vccd1 _5084_/X sky130_fd_sc_hd__o31a_1
X_8912_ _8912_/A _4436_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[21] sky130_fd_sc_hd__ebufn_8
X_8843_ _8843_/A _4355_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[22] sky130_fd_sc_hd__ebufn_8
XFILLER_24_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5986_ _5986_/A _6185_/B vssd1 vssd1 vccd1 vccd1 _6277_/B sky130_fd_sc_hd__xor2_2
XFILLER_24_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7725_ _7884_/A _8125_/A vssd1 vssd1 vccd1 vccd1 _8116_/B sky130_fd_sc_hd__nand2_2
XFILLER_12_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4937_ _5231_/B _5122_/B _4937_/C vssd1 vssd1 vccd1 vccd1 _4969_/C sky130_fd_sc_hd__or3_1
XFILLER_24_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7656_ _7643_/A _7643_/B _7641_/B _7639_/X vssd1 vssd1 vccd1 vccd1 _7660_/A sky130_fd_sc_hd__a31o_2
X_4868_ _5120_/A _5193_/A vssd1 vssd1 vccd1 vccd1 _5030_/C sky130_fd_sc_hd__or2_1
XFILLER_20_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6607_ _6710_/A _6712_/A _6710_/B _6605_/X _6778_/B vssd1 vssd1 vccd1 vccd1 _6837_/B
+ sky130_fd_sc_hd__a311o_1
XFILLER_20_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7587_ _7587_/A _8707_/Q vssd1 vssd1 vccd1 vccd1 _7588_/B sky130_fd_sc_hd__or2b_1
XFILLER_4_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4799_ _5607_/B _4831_/B _4810_/A _8602_/Q vssd1 vssd1 vccd1 vccd1 _4857_/B sky130_fd_sc_hd__or4_4
XFILLER_21_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6538_ _6539_/A _8687_/Q vssd1 vssd1 vccd1 vccd1 _6545_/B sky130_fd_sc_hd__nand2_1
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6469_ _6469_/A vssd1 vssd1 vccd1 vccd1 _8685_/D sky130_fd_sc_hd__clkbuf_1
X_8208_ _8321_/A _8230_/B _8319_/C vssd1 vssd1 vccd1 vccd1 _8475_/A sky130_fd_sc_hd__o21ba_1
X_8139_ _8191_/A _8191_/B vssd1 vssd1 vccd1 vccd1 _8163_/A sky130_fd_sc_hd__xor2_1
XFILLER_87_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5840_ _5920_/A _5840_/B vssd1 vssd1 vccd1 vccd1 _5842_/B sky130_fd_sc_hd__xor2_1
XFILLER_61_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5771_ _5771_/A _5784_/B vssd1 vssd1 vccd1 vccd1 _6032_/A sky130_fd_sc_hd__xnor2_1
X_8490_ _8490_/A _8490_/B _8490_/C vssd1 vssd1 vccd1 vccd1 _8490_/X sky130_fd_sc_hd__and3_1
X_7510_ _7503_/X _8698_/Q _7498_/Y _7509_/Y vssd1 vssd1 vccd1 vccd1 _8698_/D sky130_fd_sc_hd__o22a_1
X_4722_ _4720_/X _4721_/Y _4677_/X vssd1 vssd1 vccd1 vccd1 _8600_/D sky130_fd_sc_hd__o21a_1
X_7441_ _7443_/A _7443_/B _7440_/X vssd1 vssd1 vccd1 vccd1 _7442_/B sky130_fd_sc_hd__a21oi_2
X_4653_ _4784_/A _4653_/B vssd1 vssd1 vccd1 vccd1 _8591_/D sky130_fd_sc_hd__nor2_1
X_7372_ _7398_/A _7398_/B _7399_/B vssd1 vssd1 vccd1 vccd1 _7375_/A sky130_fd_sc_hd__or3_1
X_4584_ _4648_/A _8591_/Q vssd1 vssd1 vccd1 vccd1 _4607_/A sky130_fd_sc_hd__nor2_1
X_6323_ _6323_/A _6323_/B _6323_/C _6323_/D vssd1 vssd1 vccd1 vccd1 _6323_/X sky130_fd_sc_hd__and4_1
X_6254_ _6254_/A _6254_/B vssd1 vssd1 vccd1 vccd1 _6261_/A sky130_fd_sc_hd__xor2_1
XFILLER_103_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5205_ _5201_/X _5202_/X _5204_/X vssd1 vssd1 vccd1 vccd1 _5205_/Y sky130_fd_sc_hd__o21ai_1
X_6185_ _6185_/A _6185_/B vssd1 vssd1 vccd1 vccd1 _6281_/B sky130_fd_sc_hd__xnor2_1
XFILLER_69_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5136_ _5132_/X _5134_/X _5135_/X _4881_/X _4686_/A vssd1 vssd1 vccd1 vccd1 _5136_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_29_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5067_ _4661_/A _5062_/X _5066_/Y vssd1 vssd1 vccd1 vccd1 _5067_/X sky130_fd_sc_hd__a21o_1
XFILLER_72_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8826_ _8826_/A _4333_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[5] sky130_fd_sc_hd__ebufn_8
XFILLER_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5969_ _5969_/A _5969_/B vssd1 vssd1 vccd1 vccd1 _5970_/B sky130_fd_sc_hd__xnor2_1
XFILLER_16_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7708_ _8533_/A _7708_/B vssd1 vssd1 vccd1 vccd1 _7714_/B sky130_fd_sc_hd__nand2_1
XFILLER_52_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8688_ input3/X _8688_/D vssd1 vssd1 vccd1 vccd1 _8688_/Q sky130_fd_sc_hd__dfxtp_1
X_7639_ _7604_/A _8608_/Q vssd1 vssd1 vccd1 vccd1 _7639_/X sky130_fd_sc_hd__and2b_1
XFILLER_20_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8747__25 vssd1 vssd1 vccd1 vccd1 _8747__25/HI _8842_/A sky130_fd_sc_hd__conb_1
XFILLER_75_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7990_ _8166_/A _8063_/A vssd1 vssd1 vccd1 vccd1 _7996_/A sky130_fd_sc_hd__xor2_2
XFILLER_26_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6941_ _6938_/Y _6939_/X _6896_/X _6897_/Y vssd1 vssd1 vccd1 vccd1 _6964_/B sky130_fd_sc_hd__o211a_1
XFILLER_19_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6872_ _7137_/B _6872_/B vssd1 vssd1 vccd1 vccd1 _6876_/C sky130_fd_sc_hd__or2_1
XFILLER_62_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5823_ _5867_/A _5867_/B vssd1 vssd1 vccd1 vccd1 _5844_/A sky130_fd_sc_hd__xor2_1
XFILLER_34_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8611_ input3/X _8611_/D vssd1 vssd1 vccd1 vccd1 _8611_/Q sky130_fd_sc_hd__dfxtp_1
X_8542_ _8542_/A _8542_/B vssd1 vssd1 vccd1 vccd1 _8542_/X sky130_fd_sc_hd__xor2_1
XFILLER_22_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5754_ _5754_/A _5754_/B vssd1 vssd1 vccd1 vccd1 _5755_/D sky130_fd_sc_hd__or2_1
X_8473_ _8473_/A _8473_/B vssd1 vssd1 vccd1 vccd1 _8480_/A sky130_fd_sc_hd__xnor2_1
X_5685_ _6180_/A _5755_/B _5675_/B vssd1 vssd1 vccd1 vccd1 _5685_/Y sky130_fd_sc_hd__o21ai_1
X_4705_ _4705_/A _4994_/A vssd1 vssd1 vccd1 vccd1 _5127_/B sky130_fd_sc_hd__nor2_1
X_7424_ _7424_/A _7424_/B vssd1 vssd1 vccd1 vccd1 _7431_/B sky130_fd_sc_hd__xnor2_1
X_4636_ _8587_/Q _4637_/C _4635_/Y vssd1 vssd1 vccd1 vccd1 _8587_/D sky130_fd_sc_hd__a21oi_1
X_7355_ _7355_/A _7360_/B vssd1 vssd1 vccd1 vccd1 _7357_/B sky130_fd_sc_hd__xnor2_1
X_4567_ _8619_/Q _4567_/B vssd1 vssd1 vccd1 vccd1 _4568_/A sky130_fd_sc_hd__and2_1
X_6306_ _6306_/A _6306_/B vssd1 vssd1 vccd1 vccd1 _6326_/A sky130_fd_sc_hd__xor2_2
X_7286_ _7287_/A _7287_/B vssd1 vssd1 vccd1 vccd1 _7488_/A sky130_fd_sc_hd__nor2_1
XFILLER_89_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4498_ _7908_/B vssd1 vssd1 vccd1 vccd1 _4782_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6237_ _6237_/A _6237_/B vssd1 vssd1 vccd1 vccd1 _6238_/B sky130_fd_sc_hd__xor2_1
XFILLER_103_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6168_ _6307_/A _6106_/A _6307_/B vssd1 vssd1 vccd1 vccd1 _6168_/X sky130_fd_sc_hd__o21a_1
XFILLER_94_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5119_ _5119_/A _5119_/B _5119_/C vssd1 vssd1 vccd1 vccd1 _5120_/D sky130_fd_sc_hd__or3_1
XFILLER_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6099_ _6099_/A _6099_/B vssd1 vssd1 vccd1 vccd1 _6099_/Y sky130_fd_sc_hd__nand2_1
XFILLER_72_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5470_ _6357_/A _7699_/B _6560_/B _6351_/A vssd1 vssd1 vccd1 vccd1 _5470_/X sky130_fd_sc_hd__o211a_1
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4421_ _4427_/A vssd1 vssd1 vccd1 vccd1 _4426_/A sky130_fd_sc_hd__buf_4
XFILLER_98_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4352_ _4352_/A vssd1 vssd1 vccd1 vccd1 _4352_/Y sky130_fd_sc_hd__inv_2
X_7140_ _7140_/A _7140_/B vssd1 vssd1 vccd1 vccd1 _7141_/B sky130_fd_sc_hd__xnor2_1
XFILLER_98_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7071_ _6932_/A _6932_/B _6932_/C _6931_/B _6931_/A vssd1 vssd1 vccd1 vccd1 _7072_/C
+ sky130_fd_sc_hd__a32o_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6022_ _6199_/A _6199_/B vssd1 vssd1 vccd1 vccd1 _6023_/B sky130_fd_sc_hd__xor2_1
XFILLER_67_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7973_ _8134_/B _7973_/B vssd1 vssd1 vccd1 vccd1 _8043_/B sky130_fd_sc_hd__xnor2_1
XFILLER_54_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6924_ _6814_/A _7045_/B _6689_/A _7293_/B vssd1 vssd1 vccd1 vccd1 _6925_/C sky130_fd_sc_hd__a2bb2o_1
XFILLER_54_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6855_ _7265_/B _7092_/C vssd1 vssd1 vccd1 vccd1 _7088_/B sky130_fd_sc_hd__or2_1
XFILLER_50_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6786_ _6878_/A _6878_/B vssd1 vssd1 vccd1 vccd1 _6787_/B sky130_fd_sc_hd__xor2_1
X_5806_ _5889_/B _5890_/B vssd1 vssd1 vccd1 vccd1 _5814_/A sky130_fd_sc_hd__xnor2_1
X_8525_ _7503_/X _8717_/Q _8514_/X _8524_/X vssd1 vssd1 vccd1 vccd1 _8717_/D sky130_fd_sc_hd__o22a_1
X_5737_ _5820_/B _5737_/B vssd1 vssd1 vccd1 vccd1 _5738_/B sky130_fd_sc_hd__nand2_1
XFILLER_22_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8456_ _8417_/A _8417_/B _8416_/A vssd1 vssd1 vccd1 vccd1 _8466_/A sky130_fd_sc_hd__a21oi_1
XFILLER_13_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7407_ _7416_/B _7416_/A vssd1 vssd1 vccd1 vccd1 _7409_/B sky130_fd_sc_hd__and2b_1
X_5668_ _5754_/B _6110_/B _5706_/A _6063_/A vssd1 vssd1 vccd1 vccd1 _5675_/A sky130_fd_sc_hd__a31o_1
X_8387_ _8388_/A _8388_/B _8388_/C vssd1 vssd1 vccd1 vccd1 _8389_/A sky130_fd_sc_hd__a21oi_1
X_5599_ _5599_/A _5599_/B vssd1 vssd1 vccd1 vccd1 _5600_/B sky130_fd_sc_hd__nor2_1
X_4619_ _8582_/Q _8581_/Q _4619_/C vssd1 vssd1 vccd1 vccd1 _4623_/B sky130_fd_sc_hd__and3_1
X_7338_ _7337_/C _7337_/B _7330_/A vssd1 vssd1 vccd1 vccd1 _7345_/B sky130_fd_sc_hd__a21boi_1
X_7269_ _7268_/B _7268_/C _7268_/A vssd1 vssd1 vccd1 vccd1 _7336_/D sky130_fd_sc_hd__a21oi_1
X_8727__5 vssd1 vssd1 vccd1 vccd1 _8727__5/HI _8822_/A sky130_fd_sc_hd__conb_1
XFILLER_89_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4970_ _4970_/A _5219_/B _4970_/C _4987_/C vssd1 vssd1 vccd1 vccd1 _4970_/X sky130_fd_sc_hd__or4_1
XFILLER_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6640_ _6947_/A vssd1 vssd1 vccd1 vccd1 _7020_/A sky130_fd_sc_hd__buf_2
XFILLER_32_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6571_ _6591_/A _6580_/B vssd1 vssd1 vccd1 vccd1 _7165_/A sky130_fd_sc_hd__xor2_1
XFILLER_32_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8310_ _8310_/A _8310_/B vssd1 vssd1 vccd1 vccd1 _8379_/B sky130_fd_sc_hd__xnor2_2
X_5522_ _5794_/B _5794_/C vssd1 vssd1 vccd1 vccd1 _6006_/A sky130_fd_sc_hd__nand2_1
X_8241_ _8241_/A _8241_/B vssd1 vssd1 vccd1 vccd1 _8272_/B sky130_fd_sc_hd__xnor2_1
X_5453_ _8595_/Q _8658_/Q vssd1 vssd1 vccd1 vccd1 _5584_/A sky130_fd_sc_hd__nand2b_4
X_8172_ _8172_/A _8172_/B _8172_/C vssd1 vssd1 vccd1 vccd1 _8172_/Y sky130_fd_sc_hd__nor3_1
X_4404_ _4408_/A vssd1 vssd1 vccd1 vccd1 _4404_/Y sky130_fd_sc_hd__inv_2
X_5384_ _6357_/A _6364_/B vssd1 vssd1 vccd1 vccd1 _5384_/Y sky130_fd_sc_hd__nand2_1
XFILLER_99_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7123_ _7123_/A _7123_/B vssd1 vssd1 vccd1 vccd1 _7123_/Y sky130_fd_sc_hd__xnor2_1
X_4335_ _4339_/A vssd1 vssd1 vccd1 vccd1 _4335_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7054_ _6925_/B _6925_/C _6925_/A vssd1 vssd1 vccd1 vccd1 _7055_/C sky130_fd_sc_hd__a21bo_1
XFILLER_39_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6005_ _6005_/A _6005_/B vssd1 vssd1 vccd1 vccd1 _6224_/A sky130_fd_sc_hd__nor2_2
X_8801__79 vssd1 vssd1 vccd1 vccd1 _8801__79/HI _8910_/A sky130_fd_sc_hd__conb_1
XFILLER_27_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7956_ _8209_/A _8111_/B _8111_/C _7856_/A _7764_/A vssd1 vssd1 vccd1 vccd1 _7958_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_82_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7887_ _7887_/A _8115_/A vssd1 vssd1 vccd1 vccd1 _7963_/A sky130_fd_sc_hd__or2_1
X_6907_ _7045_/A _6907_/B _6907_/C vssd1 vssd1 vccd1 vccd1 _7057_/A sky130_fd_sc_hd__nand3b_1
XFILLER_23_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6838_ _6837_/A _6837_/B _6837_/C vssd1 vssd1 vccd1 vccd1 _6839_/B sky130_fd_sc_hd__a21o_1
XFILLER_50_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6769_ _6769_/A _6769_/B _6769_/C vssd1 vssd1 vccd1 vccd1 _6769_/X sky130_fd_sc_hd__and3_1
X_8508_ _8508_/A _8508_/B vssd1 vssd1 vccd1 vccd1 _8508_/X sky130_fd_sc_hd__xor2_1
X_8439_ _8439_/A _8439_/B vssd1 vssd1 vccd1 vccd1 _8488_/A sky130_fd_sc_hd__xnor2_1
XFILLER_2_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7810_ _7942_/A _7810_/B vssd1 vssd1 vccd1 vccd1 _7812_/B sky130_fd_sc_hd__nand2_1
XFILLER_64_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7741_ _7862_/A _8125_/A vssd1 vssd1 vccd1 vccd1 _7741_/Y sky130_fd_sc_hd__nand2_1
X_4953_ _4953_/A vssd1 vssd1 vccd1 vccd1 _4953_/X sky130_fd_sc_hd__clkbuf_2
X_7672_ _7816_/B _7666_/C _7666_/A vssd1 vssd1 vccd1 vccd1 _7687_/B sky130_fd_sc_hd__o21a_1
X_6623_ _8609_/Q _8692_/Q vssd1 vssd1 vccd1 vccd1 _6624_/B sky130_fd_sc_hd__or2b_1
X_4884_ _5068_/A vssd1 vssd1 vccd1 vccd1 _5194_/A sky130_fd_sc_hd__clkbuf_2
X_6554_ _6592_/A _6592_/B vssd1 vssd1 vccd1 vccd1 _6744_/A sky130_fd_sc_hd__nand2_2
XFILLER_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6485_ _6711_/A _7525_/A vssd1 vssd1 vccd1 vccd1 _7526_/A sky130_fd_sc_hd__or2b_1
X_5505_ _5549_/A _8601_/Q vssd1 vssd1 vccd1 vccd1 _5506_/B sky130_fd_sc_hd__nor2_1
X_8224_ _8224_/A _8224_/B vssd1 vssd1 vccd1 vccd1 _8236_/A sky130_fd_sc_hd__xnor2_1
XFILLER_10_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5436_ _5442_/A _5437_/B _5437_/C vssd1 vssd1 vccd1 vccd1 _5436_/X sky130_fd_sc_hd__a21o_1
X_8155_ _8155_/A _8383_/A vssd1 vssd1 vccd1 vccd1 _8156_/B sky130_fd_sc_hd__or2_1
XFILLER_87_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5367_ _8640_/Q _5365_/A _5357_/X vssd1 vssd1 vccd1 vccd1 _5368_/B sky130_fd_sc_hd__o21ai_1
X_8086_ _8086_/A _8086_/B vssd1 vssd1 vccd1 vccd1 _8087_/B sky130_fd_sc_hd__nand2_1
X_5298_ _8622_/Q _5300_/B vssd1 vssd1 vccd1 vccd1 _5298_/X sky130_fd_sc_hd__or2_1
X_7106_ _7106_/A _7106_/B vssd1 vssd1 vccd1 vccd1 _7112_/A sky130_fd_sc_hd__xnor2_1
XFILLER_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7037_ _7037_/A _7129_/B vssd1 vssd1 vccd1 vccd1 _7042_/A sky130_fd_sc_hd__xnor2_1
XFILLER_28_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7939_ _7938_/A _7938_/B _7938_/C vssd1 vssd1 vccd1 vccd1 _7940_/B sky130_fd_sc_hd__o21a_1
XFILLER_15_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6270_ _6270_/A _6270_/B vssd1 vssd1 vccd1 vccd1 _6271_/B sky130_fd_sc_hd__xnor2_1
XFILLER_103_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5221_ _4970_/A _5218_/X _5220_/X vssd1 vssd1 vccd1 vccd1 _5221_/X sky130_fd_sc_hd__o21a_1
X_5152_ _5190_/B _5152_/B _5163_/A vssd1 vssd1 vccd1 vccd1 _5152_/Y sky130_fd_sc_hd__nor3b_2
XFILLER_96_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5083_ _5083_/A _5231_/B _5120_/A _5166_/B vssd1 vssd1 vccd1 vccd1 _5083_/X sky130_fd_sc_hd__or4_1
X_8911_ _8911_/A _4435_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[20] sky130_fd_sc_hd__ebufn_8
X_8842_ _8842_/A _4354_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[21] sky130_fd_sc_hd__ebufn_8
XFILLER_37_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7724_ _7862_/B vssd1 vssd1 vccd1 vccd1 _8125_/A sky130_fd_sc_hd__clkbuf_2
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5985_ _5985_/A _6203_/B vssd1 vssd1 vccd1 vccd1 _6185_/B sky130_fd_sc_hd__and2_1
XFILLER_40_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4936_ _5041_/A _4955_/B _5230_/B vssd1 vssd1 vccd1 vccd1 _5122_/B sky130_fd_sc_hd__o21ai_2
X_7655_ _7988_/A vssd1 vssd1 vccd1 vccd1 _7671_/A sky130_fd_sc_hd__clkbuf_2
X_4867_ _5241_/B _5231_/C vssd1 vssd1 vccd1 vccd1 _5193_/A sky130_fd_sc_hd__or2_2
XFILLER_20_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6606_ _7529_/A _7688_/B vssd1 vssd1 vccd1 vccd1 _6778_/B sky130_fd_sc_hd__nor2_1
X_7586_ _8707_/Q _7587_/A vssd1 vssd1 vccd1 vccd1 _7588_/A sky130_fd_sc_hd__or2b_1
X_4798_ _4752_/A _4903_/A _4897_/C vssd1 vssd1 vccd1 vccd1 _4916_/B sky130_fd_sc_hd__a21oi_4
X_6537_ _6513_/A _6545_/A _6534_/X _6536_/X vssd1 vssd1 vccd1 vccd1 _8692_/D sky130_fd_sc_hd__a31o_1
X_6468_ _6466_/Y _6468_/B vssd1 vssd1 vccd1 vccd1 _6469_/A sky130_fd_sc_hd__and2b_1
X_8207_ _8207_/A _8230_/B vssd1 vssd1 vccd1 vccd1 _8319_/C sky130_fd_sc_hd__and2_1
X_5419_ _5419_/A vssd1 vssd1 vccd1 vccd1 _5419_/X sky130_fd_sc_hd__clkbuf_2
X_6399_ _8684_/Q _6399_/B _8685_/Q _8683_/Q vssd1 vssd1 vccd1 vccd1 _6400_/C sky130_fd_sc_hd__and4b_1
X_8138_ _8138_/A _8138_/B vssd1 vssd1 vccd1 vccd1 _8191_/B sky130_fd_sc_hd__xnor2_2
XFILLER_101_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8069_ _8069_/A _8069_/B vssd1 vssd1 vccd1 vccd1 _8070_/B sky130_fd_sc_hd__or2_1
XFILLER_75_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5770_ _5770_/A _5770_/B vssd1 vssd1 vccd1 vccd1 _5784_/B sky130_fd_sc_hd__xor2_1
X_4721_ _5265_/A _4724_/S vssd1 vssd1 vccd1 vccd1 _4721_/Y sky130_fd_sc_hd__nor2_1
X_7440_ _7439_/A _7440_/B vssd1 vssd1 vccd1 vccd1 _7440_/X sky130_fd_sc_hd__and2b_1
X_4652_ _8591_/Q _4646_/C _5402_/C vssd1 vssd1 vccd1 vccd1 _4653_/B sky130_fd_sc_hd__o21a_1
X_7371_ _7378_/D _7371_/B vssd1 vssd1 vccd1 vccd1 _7399_/B sky130_fd_sc_hd__xnor2_1
X_4583_ input2/X vssd1 vssd1 vccd1 vccd1 _4648_/A sky130_fd_sc_hd__inv_2
X_6322_ _6322_/A _6322_/B vssd1 vssd1 vccd1 vccd1 _6322_/X sky130_fd_sc_hd__or2_1
X_6253_ _6215_/A _6215_/B _6215_/C _6218_/B _6218_/A vssd1 vssd1 vccd1 vccd1 _6254_/B
+ sky130_fd_sc_hd__o32a_1
XFILLER_88_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5204_ _5166_/D _5168_/X _5203_/Y _4731_/A _5185_/A vssd1 vssd1 vccd1 vccd1 _5204_/X
+ sky130_fd_sc_hd__o221a_1
X_6184_ _6183_/Y _5982_/B _5980_/X vssd1 vssd1 vccd1 vccd1 _6186_/A sky130_fd_sc_hd__a21boi_1
X_5135_ _5135_/A _5166_/A _5135_/C _5135_/D vssd1 vssd1 vccd1 vccd1 _5135_/X sky130_fd_sc_hd__or4_1
XFILLER_57_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5066_ _5066_/A _5066_/B vssd1 vssd1 vccd1 vccd1 _5066_/Y sky130_fd_sc_hd__nand2_1
XFILLER_44_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8825_ _8825_/A _4332_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[4] sky130_fd_sc_hd__ebufn_8
XFILLER_80_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5968_ _6180_/B _5968_/B vssd1 vssd1 vccd1 vccd1 _5969_/B sky130_fd_sc_hd__xnor2_1
XFILLER_40_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7707_ _8719_/Q vssd1 vssd1 vccd1 vccd1 _8533_/A sky130_fd_sc_hd__inv_2
X_4919_ _5180_/C vssd1 vssd1 vccd1 vccd1 _5137_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_40_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8687_ input3/X _8687_/D vssd1 vssd1 vccd1 vccd1 _8687_/Q sky130_fd_sc_hd__dfxtp_1
X_5899_ _5900_/A _5900_/B _5900_/C vssd1 vssd1 vccd1 vccd1 _5901_/A sky130_fd_sc_hd__o21a_1
X_7638_ _7649_/A _7654_/B _7633_/X _7631_/X vssd1 vssd1 vccd1 vccd1 _7643_/B sky130_fd_sc_hd__a211o_1
XFILLER_20_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7569_ _8711_/Q vssd1 vssd1 vccd1 vccd1 _7604_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_79_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6940_ _6896_/X _6897_/Y _6938_/Y _6939_/X vssd1 vssd1 vccd1 vccd1 _6964_/A sky130_fd_sc_hd__a211oi_2
XFILLER_93_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6871_ _7174_/B _7197_/B _6870_/X vssd1 vssd1 vccd1 vccd1 _6872_/B sky130_fd_sc_hd__a21bo_1
XFILLER_62_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8610_ input3/X _8610_/D vssd1 vssd1 vccd1 vccd1 _8610_/Q sky130_fd_sc_hd__dfxtp_1
X_5822_ _5822_/A _5822_/B vssd1 vssd1 vccd1 vccd1 _5867_/B sky130_fd_sc_hd__xnor2_2
X_8541_ _8531_/A _8539_/B _8532_/Y vssd1 vssd1 vccd1 vccd1 _8542_/B sky130_fd_sc_hd__a21o_1
X_5753_ _5753_/A _5753_/B vssd1 vssd1 vccd1 vccd1 _5755_/C sky130_fd_sc_hd__xnor2_1
X_4704_ _4705_/A _4994_/A vssd1 vssd1 vccd1 vccd1 _5127_/A sky130_fd_sc_hd__and2_1
X_8472_ _8472_/A _8472_/B vssd1 vssd1 vccd1 vccd1 _8473_/B sky130_fd_sc_hd__xnor2_1
X_5684_ _5749_/B vssd1 vssd1 vccd1 vccd1 _5755_/B sky130_fd_sc_hd__clkbuf_2
X_7423_ _7423_/A _7423_/B vssd1 vssd1 vccd1 vccd1 _7424_/B sky130_fd_sc_hd__nand2_1
X_4635_ _8587_/Q _4637_/C _4646_/A vssd1 vssd1 vccd1 vccd1 _4635_/Y sky130_fd_sc_hd__o21ai_1
X_7354_ _7354_/A _7354_/B vssd1 vssd1 vccd1 vccd1 _7360_/B sky130_fd_sc_hd__xor2_1
X_4566_ _4566_/A vssd1 vssd1 vccd1 vccd1 _8872_/A sky130_fd_sc_hd__clkbuf_1
X_6305_ _6301_/X _6337_/A _6304_/X vssd1 vssd1 vccd1 vccd1 _6320_/A sky130_fd_sc_hd__o21a_1
XFILLER_103_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7285_ _7283_/A _7283_/B _7284_/X vssd1 vssd1 vccd1 vccd1 _7287_/B sky130_fd_sc_hd__a21oi_1
X_4497_ _7783_/A vssd1 vssd1 vccd1 vccd1 _7908_/B sky130_fd_sc_hd__clkbuf_4
X_6236_ _6288_/B _6236_/B vssd1 vssd1 vccd1 vccd1 _6237_/B sky130_fd_sc_hd__xnor2_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6167_ _6167_/A vssd1 vssd1 vccd1 vccd1 _6307_/A sky130_fd_sc_hd__inv_2
XFILLER_85_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5118_ _8592_/Q _5118_/B _5118_/C _5118_/D vssd1 vssd1 vccd1 vccd1 _5118_/X sky130_fd_sc_hd__or4_1
XFILLER_72_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6098_ _6099_/A _6099_/B vssd1 vssd1 vccd1 vccd1 _6157_/B sky130_fd_sc_hd__xnor2_2
XFILLER_84_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5049_ _5057_/A _5174_/B _5165_/C _5049_/D vssd1 vssd1 vccd1 vccd1 _5049_/X sky130_fd_sc_hd__or4_1
XFILLER_38_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8807__85 vssd1 vssd1 vccd1 vccd1 _8807__85/HI _8916_/A sky130_fd_sc_hd__conb_1
XFILLER_76_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4420_ _4420_/A vssd1 vssd1 vccd1 vccd1 _4420_/Y sky130_fd_sc_hd__inv_2
X_4351_ _4352_/A vssd1 vssd1 vccd1 vccd1 _4351_/Y sky130_fd_sc_hd__inv_2
X_7070_ _7101_/D _7069_/B _7069_/C vssd1 vssd1 vccd1 vccd1 _7072_/B sky130_fd_sc_hd__a21o_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6021_ _6021_/A _6021_/B vssd1 vssd1 vccd1 vccd1 _6199_/B sky130_fd_sc_hd__xor2_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7972_ _7972_/A _7972_/B vssd1 vssd1 vccd1 vccd1 _7973_/B sky130_fd_sc_hd__xor2_1
XFILLER_27_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6923_ _7062_/B _6922_/C _6922_/A vssd1 vssd1 vccd1 vccd1 _6925_/B sky130_fd_sc_hd__a21o_1
XFILLER_35_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6854_ _6854_/A _6854_/B vssd1 vssd1 vccd1 vccd1 _7159_/A sky130_fd_sc_hd__xnor2_1
XFILLER_35_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6785_ _6785_/A _6825_/B vssd1 vssd1 vccd1 vccd1 _6878_/B sky130_fd_sc_hd__xor2_1
XFILLER_50_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5805_ _5805_/A _5805_/B vssd1 vssd1 vccd1 vccd1 _5890_/B sky130_fd_sc_hd__xnor2_1
X_8524_ _8527_/A _8527_/B _8524_/C vssd1 vssd1 vccd1 vccd1 _8524_/X sky130_fd_sc_hd__and3_1
X_5736_ _5736_/A _5736_/B vssd1 vssd1 vccd1 vccd1 _5737_/B sky130_fd_sc_hd__or2_1
X_8455_ _8455_/A _8455_/B vssd1 vssd1 vccd1 vccd1 _8481_/A sky130_fd_sc_hd__xnor2_1
X_5667_ _5961_/A vssd1 vssd1 vccd1 vccd1 _6110_/B sky130_fd_sc_hd__clkbuf_2
X_7406_ _7402_/A _7402_/B _7423_/A vssd1 vssd1 vccd1 vccd1 _7416_/A sky130_fd_sc_hd__a21bo_1
X_4618_ _8581_/Q _4619_/C _4617_/Y vssd1 vssd1 vccd1 vccd1 _8581_/D sky130_fd_sc_hd__a21oi_1
X_8386_ _8472_/A _8386_/B vssd1 vssd1 vccd1 vccd1 _8388_/C sky130_fd_sc_hd__nor2_1
X_5598_ _5740_/A _5740_/B vssd1 vssd1 vccd1 vccd1 _5599_/B sky130_fd_sc_hd__nor2_1
X_4549_ _4549_/A vssd1 vssd1 vccd1 vccd1 _8868_/A sky130_fd_sc_hd__clkbuf_1
X_7337_ _7330_/A _7337_/B _7337_/C vssd1 vssd1 vccd1 vccd1 _7345_/A sky130_fd_sc_hd__and3b_1
XFILLER_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7268_ _7268_/A _7268_/B _7268_/C vssd1 vssd1 vccd1 vccd1 _7336_/C sky130_fd_sc_hd__and3_1
XFILLER_104_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6219_ _6249_/A _6249_/B vssd1 vssd1 vccd1 vccd1 _6222_/A sky130_fd_sc_hd__xnor2_2
X_7199_ _7226_/B _7199_/B vssd1 vssd1 vccd1 vccd1 _7234_/B sky130_fd_sc_hd__and2_1
XFILLER_58_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_10 _7676_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6570_ _8689_/Q _8606_/Q vssd1 vssd1 vccd1 vccd1 _6580_/B sky130_fd_sc_hd__xnor2_4
XFILLER_32_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5521_ _5580_/B vssd1 vssd1 vccd1 vccd1 _6005_/A sky130_fd_sc_hd__clkbuf_2
X_8240_ _8240_/A _8299_/B vssd1 vssd1 vccd1 vccd1 _8241_/B sky130_fd_sc_hd__xnor2_1
X_5452_ _5452_/A vssd1 vssd1 vccd1 vccd1 _8653_/D sky130_fd_sc_hd__clkbuf_1
X_8171_ _8382_/A _8196_/A vssd1 vssd1 vccd1 vccd1 _8172_/C sky130_fd_sc_hd__nor2_1
X_4403_ _4427_/A vssd1 vssd1 vccd1 vccd1 _4408_/A sky130_fd_sc_hd__buf_6
X_5383_ _8645_/Q vssd1 vssd1 vccd1 vccd1 _6364_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_7122_ _7306_/A _7122_/B vssd1 vssd1 vccd1 vccd1 _7123_/B sky130_fd_sc_hd__xnor2_1
X_4334_ _4459_/A vssd1 vssd1 vccd1 vccd1 _4339_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_99_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7053_ _7051_/B _7051_/C _7099_/A vssd1 vssd1 vccd1 vccd1 _7101_/B sky130_fd_sc_hd__o21ai_2
XFILLER_5_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6004_ _5896_/A _5540_/B _6226_/A _5587_/Y vssd1 vssd1 vccd1 vccd1 _6008_/A sky130_fd_sc_hd__a31o_1
XFILLER_101_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8798__76 vssd1 vssd1 vccd1 vccd1 _8798__76/HI _8907_/A sky130_fd_sc_hd__conb_1
XFILLER_67_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7955_ _7972_/B vssd1 vssd1 vccd1 vccd1 _8117_/S sky130_fd_sc_hd__clkbuf_2
X_7886_ _7886_/A _7962_/B _7886_/C vssd1 vssd1 vccd1 vccd1 _7892_/B sky130_fd_sc_hd__and3_1
X_6906_ _6905_/B _6905_/C _7045_/B vssd1 vssd1 vccd1 vccd1 _6907_/C sky130_fd_sc_hd__o21ai_1
XFILLER_35_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6837_ _6837_/A _6837_/B _6837_/C vssd1 vssd1 vccd1 vccd1 _6839_/A sky130_fd_sc_hd__nand3_1
X_8507_ _8489_/Y _8490_/X _8494_/X _8506_/X vssd1 vssd1 vccd1 vccd1 _8527_/B sky130_fd_sc_hd__o211a_2
X_6768_ _6769_/C _6768_/B vssd1 vssd1 vccd1 vccd1 _6768_/X sky130_fd_sc_hd__and2b_1
X_6699_ _6724_/A _6703_/C _7180_/A vssd1 vssd1 vccd1 vccd1 _7163_/B sky130_fd_sc_hd__a21o_1
X_5719_ _5717_/X _5601_/B _5718_/Y vssd1 vssd1 vccd1 vccd1 _5739_/A sky130_fd_sc_hd__a21boi_2
X_8438_ _8438_/A _8438_/B vssd1 vssd1 vccd1 vccd1 _8439_/B sky130_fd_sc_hd__xnor2_1
X_8369_ _8290_/A _8290_/B _8368_/X vssd1 vssd1 vccd1 vccd1 _8370_/B sky130_fd_sc_hd__a21oi_1
XFILLER_49_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7740_ _7740_/A _7740_/B vssd1 vssd1 vccd1 vccd1 _7862_/A sky130_fd_sc_hd__xnor2_2
X_4952_ _4952_/A _5113_/A vssd1 vssd1 vccd1 vccd1 _4953_/A sky130_fd_sc_hd__nor2_1
X_7671_ _7671_/A vssd1 vssd1 vccd1 vccd1 _7816_/B sky130_fd_sc_hd__clkbuf_2
X_4883_ _5240_/A vssd1 vssd1 vccd1 vccd1 _5075_/B sky130_fd_sc_hd__buf_2
XFILLER_32_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6622_ _8692_/Q _8609_/Q vssd1 vssd1 vccd1 vccd1 _6626_/A sky130_fd_sc_hd__or2b_1
XFILLER_20_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6553_ _7511_/S _7708_/B vssd1 vssd1 vccd1 vccd1 _6592_/B sky130_fd_sc_hd__nand2_1
XFILLER_9_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6484_ _8702_/Q vssd1 vssd1 vccd1 vccd1 _6711_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5504_ _5549_/A _8601_/Q vssd1 vssd1 vccd1 vccd1 _5506_/A sky130_fd_sc_hd__and2_1
X_8223_ _8315_/A _8315_/B vssd1 vssd1 vccd1 vccd1 _8224_/B sky130_fd_sc_hd__xnor2_1
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5435_ _5428_/A _5433_/B _5434_/X vssd1 vssd1 vccd1 vccd1 _5437_/C sky130_fd_sc_hd__o21a_1
X_8154_ _8155_/A _8383_/A vssd1 vssd1 vccd1 vccd1 _8202_/A sky130_fd_sc_hd__nand2_1
XFILLER_59_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5366_ _8639_/Q _8640_/Q _5366_/C vssd1 vssd1 vccd1 vccd1 _5369_/B sky130_fd_sc_hd__and3_1
X_8085_ _8086_/A _8086_/B vssd1 vssd1 vccd1 vccd1 _8185_/A sky130_fd_sc_hd__or2_1
X_5297_ _8696_/Q _5285_/X _5295_/X _5296_/X vssd1 vssd1 vccd1 vccd1 _8621_/D sky130_fd_sc_hd__o211a_1
X_7105_ _7105_/A _7105_/B vssd1 vssd1 vccd1 vccd1 _7106_/B sky130_fd_sc_hd__xnor2_1
XFILLER_87_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7036_ _7036_/A _7036_/B vssd1 vssd1 vccd1 vccd1 _7129_/B sky130_fd_sc_hd__xnor2_1
XFILLER_28_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7938_ _7938_/A _7938_/B _7938_/C vssd1 vssd1 vccd1 vccd1 _7940_/A sky130_fd_sc_hd__nor3_1
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7869_ _7869_/A _7869_/B vssd1 vssd1 vccd1 vccd1 _8326_/A sky130_fd_sc_hd__xnor2_2
XFILLER_11_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5220_ _5070_/D _5219_/X _5074_/X vssd1 vssd1 vccd1 vccd1 _5220_/X sky130_fd_sc_hd__a21o_1
XFILLER_102_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5151_ _5151_/A _5151_/B _5180_/C vssd1 vssd1 vccd1 vccd1 _5163_/A sky130_fd_sc_hd__nor3_1
XFILLER_69_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5082_ _5067_/X _5070_/X _5073_/X _5081_/X vssd1 vssd1 vccd1 vccd1 _5082_/X sky130_fd_sc_hd__a31o_1
XFILLER_96_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8910_ _8910_/A _4434_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[19] sky130_fd_sc_hd__ebufn_8
XFILLER_77_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8768__46 vssd1 vssd1 vccd1 vccd1 _8768__46/HI _8863_/A sky130_fd_sc_hd__conb_1
XFILLER_37_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8841_ _8841_/A _4352_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[20] sky130_fd_sc_hd__ebufn_8
XFILLER_52_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7723_ _7954_/A vssd1 vssd1 vccd1 vccd1 _8134_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_52_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5984_ _5984_/A _6183_/A vssd1 vssd1 vccd1 vccd1 _6203_/B sky130_fd_sc_hd__nand2_1
X_4935_ _5015_/A _5245_/C vssd1 vssd1 vccd1 vccd1 _5230_/B sky130_fd_sc_hd__nor2_1
X_7654_ _7673_/A _7654_/B vssd1 vssd1 vccd1 vccd1 _7988_/A sky130_fd_sc_hd__xnor2_2
X_4866_ _4866_/A _4990_/B vssd1 vssd1 vccd1 vccd1 _5231_/C sky130_fd_sc_hd__nand2_2
XFILLER_20_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6605_ _8702_/Q _6605_/B vssd1 vssd1 vccd1 vccd1 _6605_/X sky130_fd_sc_hd__and2b_1
X_7585_ _7627_/A _7581_/X _7584_/Y vssd1 vssd1 vccd1 vccd1 _8708_/D sky130_fd_sc_hd__o21a_1
X_4797_ _4961_/B vssd1 vssd1 vccd1 vccd1 _4897_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_21_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6536_ _6536_/A _6536_/B _7540_/A vssd1 vssd1 vccd1 vccd1 _6536_/X sky130_fd_sc_hd__and3_1
XFILLER_97_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6467_ _8684_/Q _6465_/A _6466_/Y _4743_/X vssd1 vssd1 vccd1 vccd1 _8684_/D sky130_fd_sc_hd__o211a_1
X_8206_ _8206_/A _8462_/A vssd1 vssd1 vccd1 vccd1 _8230_/B sky130_fd_sc_hd__nor2_1
X_5418_ _5414_/A _5412_/X _5413_/X _5417_/X vssd1 vssd1 vccd1 vccd1 _8648_/D sky130_fd_sc_hd__a22o_1
X_6398_ _6398_/A _6398_/B _6398_/C vssd1 vssd1 vccd1 vccd1 _6399_/B sky130_fd_sc_hd__and3_1
XFILLER_102_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8137_ _8398_/A _8194_/B vssd1 vssd1 vccd1 vccd1 _8138_/B sky130_fd_sc_hd__xnor2_2
XFILLER_87_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5349_ _8635_/Q vssd1 vssd1 vccd1 vccd1 _6471_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_101_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8068_ _8068_/A _8068_/B vssd1 vssd1 vccd1 vccd1 _8070_/A sky130_fd_sc_hd__nand2_1
XFILLER_47_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7019_ _6914_/B _6914_/C _6914_/A vssd1 vssd1 vccd1 vccd1 _7037_/A sky130_fd_sc_hd__a21boi_1
XFILLER_46_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8782__60 vssd1 vssd1 vccd1 vccd1 _8782__60/HI _8891_/A sky130_fd_sc_hd__conb_1
XFILLER_43_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4720_ _5265_/A _4724_/S vssd1 vssd1 vccd1 vccd1 _4720_/X sky130_fd_sc_hd__and2_1
XFILLER_42_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4651_ _5406_/B vssd1 vssd1 vccd1 vccd1 _5402_/C sky130_fd_sc_hd__clkbuf_2
X_7370_ _7046_/A _7297_/B _7439_/A vssd1 vssd1 vccd1 vccd1 _7371_/B sky130_fd_sc_hd__a21oi_1
X_4582_ _8571_/Q _4582_/B vssd1 vssd1 vccd1 vccd1 _8571_/D sky130_fd_sc_hd__nor2_1
X_6321_ _6322_/A _6322_/B vssd1 vssd1 vccd1 vccd1 _6327_/A sky130_fd_sc_hd__nand2_1
X_6252_ _6227_/S _6228_/A _6251_/X vssd1 vssd1 vccd1 vccd1 _6254_/A sky130_fd_sc_hd__a21bo_1
XFILLER_88_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5203_ _5203_/A vssd1 vssd1 vccd1 vccd1 _5203_/Y sky130_fd_sc_hd__inv_2
X_6183_ _6183_/A vssd1 vssd1 vccd1 vccd1 _6183_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5134_ _5133_/Y _5159_/C _5105_/X vssd1 vssd1 vccd1 vccd1 _5134_/X sky130_fd_sc_hd__o21a_1
XFILLER_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5065_ _5214_/B _5149_/B _5137_/B _5017_/A vssd1 vssd1 vccd1 vccd1 _5066_/B sky130_fd_sc_hd__nor4b_1
X_8824_ _8824_/A _4331_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[3] sky130_fd_sc_hd__ebufn_8
XFILLER_16_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5967_ _5967_/A _5967_/B vssd1 vssd1 vccd1 vccd1 _5969_/A sky130_fd_sc_hd__xor2_1
XFILLER_80_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7706_ _7740_/A _7740_/B vssd1 vssd1 vccd1 vccd1 _7746_/A sky130_fd_sc_hd__xor2_2
XFILLER_12_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4918_ _4946_/A vssd1 vssd1 vccd1 vccd1 _5098_/D sky130_fd_sc_hd__clkbuf_2
X_8686_ input3/X _8686_/D vssd1 vssd1 vccd1 vccd1 _8686_/Q sky130_fd_sc_hd__dfxtp_1
X_7637_ _7779_/A vssd1 vssd1 vccd1 vccd1 _7986_/A sky130_fd_sc_hd__clkbuf_2
X_5898_ _5898_/A _5898_/B vssd1 vssd1 vccd1 vccd1 _5900_/C sky130_fd_sc_hd__xnor2_1
X_4849_ _4849_/A _4849_/B vssd1 vssd1 vccd1 vccd1 _5026_/B sky130_fd_sc_hd__nor2_1
X_7568_ _8709_/Q vssd1 vssd1 vccd1 vccd1 _7587_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7499_ _6334_/X _8695_/Q _7493_/Y _7498_/Y vssd1 vssd1 vccd1 vccd1 _8695_/D sky130_fd_sc_hd__o22a_1
X_6519_ _6520_/A _6526_/B vssd1 vssd1 vccd1 vccd1 _6521_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8738__16 vssd1 vssd1 vccd1 vccd1 _8738__16/HI _8833_/A sky130_fd_sc_hd__conb_1
X_6870_ _7223_/B _6883_/B vssd1 vssd1 vccd1 vccd1 _6870_/X sky130_fd_sc_hd__or2_1
XFILLER_81_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5821_ _5875_/A _5821_/B vssd1 vssd1 vccd1 vccd1 _5822_/B sky130_fd_sc_hd__and2_1
X_8540_ _8540_/A _8540_/B vssd1 vssd1 vccd1 vccd1 _8542_/A sky130_fd_sc_hd__nor2_1
XFILLER_62_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5752_ _5674_/A _6180_/B _5751_/X vssd1 vssd1 vccd1 vccd1 _5753_/B sky130_fd_sc_hd__o21ba_1
XFILLER_22_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4703_ _4662_/A _4697_/Y _4702_/X _4677_/X vssd1 vssd1 vccd1 vccd1 _8596_/D sky130_fd_sc_hd__o211a_1
X_8471_ _8471_/A _8471_/B vssd1 vssd1 vccd1 vccd1 _8472_/B sky130_fd_sc_hd__xnor2_1
X_5683_ _5961_/B vssd1 vssd1 vccd1 vccd1 _5749_/B sky130_fd_sc_hd__clkbuf_2
X_7422_ _7422_/A _7422_/B vssd1 vssd1 vccd1 vccd1 _7423_/B sky130_fd_sc_hd__nand2_1
X_4634_ _4637_/C _4634_/B vssd1 vssd1 vccd1 vccd1 _8586_/D sky130_fd_sc_hd__nor2_1
X_7353_ _7353_/A _7353_/B vssd1 vssd1 vccd1 vccd1 _7354_/B sky130_fd_sc_hd__xnor2_1
X_4565_ _8618_/Q _4567_/B vssd1 vssd1 vccd1 vccd1 _4566_/A sky130_fd_sc_hd__and2_1
X_6304_ _6316_/A _6304_/B _6304_/C vssd1 vssd1 vccd1 vccd1 _6304_/X sky130_fd_sc_hd__and3b_1
X_7284_ _7462_/A _7456_/B vssd1 vssd1 vccd1 vccd1 _7284_/X sky130_fd_sc_hd__and2_1
X_4496_ _8611_/Q vssd1 vssd1 vccd1 vccd1 _7783_/A sky130_fd_sc_hd__clkbuf_4
X_6235_ _6266_/A _6266_/B vssd1 vssd1 vccd1 vccd1 _6236_/B sky130_fd_sc_hd__xnor2_2
XFILLER_69_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6166_ _6316_/A _6316_/B _6312_/A _6165_/X vssd1 vssd1 vccd1 vccd1 _6310_/B sky130_fd_sc_hd__a31o_1
XFILLER_84_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5117_ _4990_/A _5231_/C _5202_/B _5115_/X _5116_/X vssd1 vssd1 vccd1 vccd1 _5117_/X
+ sky130_fd_sc_hd__o41a_1
X_6097_ _6097_/A _6097_/B vssd1 vssd1 vccd1 vccd1 _6099_/B sky130_fd_sc_hd__xor2_2
XFILLER_84_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5048_ _4969_/B _5044_/X _5047_/X vssd1 vssd1 vccd1 vccd1 _5049_/D sky130_fd_sc_hd__o21a_1
XFILLER_80_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6999_ _6999_/A _6999_/B vssd1 vssd1 vccd1 vccd1 _6999_/X sky130_fd_sc_hd__or2_1
XFILLER_43_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8752__30 vssd1 vssd1 vccd1 vccd1 _8752__30/HI _8847_/A sky130_fd_sc_hd__conb_1
XFILLER_21_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8669_ input3/X _8669_/D vssd1 vssd1 vccd1 vccd1 _8669_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4350_ _4352_/A vssd1 vssd1 vccd1 vccd1 _4350_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6020_ _6020_/A _6210_/A vssd1 vssd1 vccd1 vccd1 _6021_/B sky130_fd_sc_hd__xnor2_1
XFILLER_79_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7971_ _7877_/A _8406_/A _7879_/B _7879_/A vssd1 vssd1 vccd1 vccd1 _8043_/A sky130_fd_sc_hd__a22o_1
X_6922_ _6922_/A _7062_/B _6922_/C vssd1 vssd1 vccd1 vccd1 _6925_/A sky130_fd_sc_hd__nand3_1
X_6853_ _6854_/A _6854_/B vssd1 vssd1 vccd1 vccd1 _6853_/X sky130_fd_sc_hd__and2_1
X_5804_ _5812_/A _6220_/B _5903_/A vssd1 vssd1 vccd1 vccd1 _5805_/B sky130_fd_sc_hd__o21ai_1
X_6784_ _6886_/A _6784_/B vssd1 vssd1 vccd1 vccd1 _6825_/B sky130_fd_sc_hd__and2_1
XFILLER_22_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8523_ _8526_/S _8523_/B vssd1 vssd1 vccd1 vccd1 _8524_/C sky130_fd_sc_hd__nand2_1
X_5735_ _5736_/A _5736_/B vssd1 vssd1 vccd1 vccd1 _5820_/B sky130_fd_sc_hd__nand2_1
XFILLER_13_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8454_ _8419_/A _8452_/X _8453_/X vssd1 vssd1 vccd1 vccd1 _8455_/B sky130_fd_sc_hd__o21a_1
X_5666_ _5666_/A vssd1 vssd1 vccd1 vccd1 _5754_/B sky130_fd_sc_hd__clkbuf_2
X_7405_ _7422_/A _7422_/B vssd1 vssd1 vccd1 vccd1 _7423_/A sky130_fd_sc_hd__or2_1
X_4617_ _8581_/Q _4619_/C _4607_/X vssd1 vssd1 vccd1 vccd1 _4617_/Y sky130_fd_sc_hd__o21ai_1
X_8385_ _8385_/A _8385_/B _8445_/B vssd1 vssd1 vccd1 vccd1 _8386_/B sky130_fd_sc_hd__and3_1
X_5597_ _5740_/A _5740_/B vssd1 vssd1 vccd1 vccd1 _5599_/A sky130_fd_sc_hd__and2_1
X_7336_ _7336_/A _7336_/B _7336_/C _7336_/D vssd1 vssd1 vccd1 vccd1 _7337_/C sky130_fd_sc_hd__or4_1
XFILLER_89_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4548_ _8614_/Q _4552_/B vssd1 vssd1 vccd1 vccd1 _4549_/A sky130_fd_sc_hd__and2_2
XFILLER_104_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7267_ _7334_/D _7334_/C _7313_/B _7270_/A vssd1 vssd1 vccd1 vccd1 _7336_/B sky130_fd_sc_hd__o2bb2a_1
X_4479_ _8604_/Q vssd1 vssd1 vccd1 vccd1 _4831_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6218_ _6218_/A _6218_/B vssd1 vssd1 vccd1 vccd1 _6249_/B sky130_fd_sc_hd__xor2_2
X_7198_ _7227_/A _7196_/X _7305_/A vssd1 vssd1 vccd1 vccd1 _7234_/A sky130_fd_sc_hd__o21a_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6149_ _6138_/A _6149_/B vssd1 vssd1 vccd1 vccd1 _6153_/B sky130_fd_sc_hd__and2b_1
XFILLER_85_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5520_ _5520_/A _5520_/B vssd1 vssd1 vccd1 vccd1 _5580_/B sky130_fd_sc_hd__xnor2_2
X_5451_ _7547_/A _5451_/B _5451_/C vssd1 vssd1 vccd1 vccd1 _5452_/A sky130_fd_sc_hd__and3_1
X_8170_ _8302_/A vssd1 vssd1 vccd1 vccd1 _8382_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4402_ input1/X vssd1 vssd1 vccd1 vccd1 _4427_/A sky130_fd_sc_hd__clkbuf_2
X_5382_ _8661_/Q vssd1 vssd1 vccd1 vccd1 _6357_/A sky130_fd_sc_hd__inv_2
X_7121_ _7121_/A _7121_/B vssd1 vssd1 vccd1 vccd1 _7122_/B sky130_fd_sc_hd__xnor2_1
X_4333_ _4333_/A vssd1 vssd1 vccd1 vccd1 _4333_/Y sky130_fd_sc_hd__inv_2
X_7052_ _7052_/A vssd1 vssd1 vccd1 vccd1 _7115_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6003_ _6003_/A _6007_/A vssd1 vssd1 vccd1 vccd1 _6226_/A sky130_fd_sc_hd__or2_1
XFILLER_67_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7954_ _7954_/A _7954_/B vssd1 vssd1 vccd1 vccd1 _7972_/B sky130_fd_sc_hd__or2_1
XFILLER_54_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6905_ _7045_/B _6905_/B _6905_/C vssd1 vssd1 vccd1 vccd1 _6907_/B sky130_fd_sc_hd__or3_1
XFILLER_54_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7885_ _7885_/A _7972_/A vssd1 vssd1 vccd1 vccd1 _7892_/A sky130_fd_sc_hd__nor2_1
XFILLER_24_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6836_ _6836_/A _6836_/B vssd1 vssd1 vccd1 vccd1 _6837_/C sky130_fd_sc_hd__nand2_1
XFILLER_62_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6767_ _6767_/A _6767_/B vssd1 vssd1 vccd1 vccd1 _6771_/A sky130_fd_sc_hd__xor2_1
XFILLER_50_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8506_ _8497_/Y _8498_/X _8502_/Y _8505_/Y vssd1 vssd1 vccd1 vccd1 _8506_/X sky130_fd_sc_hd__o211a_1
X_5718_ _5718_/A _5718_/B vssd1 vssd1 vccd1 vccd1 _5718_/Y sky130_fd_sc_hd__nand2_1
X_6698_ _7165_/A _6723_/A _7167_/B _6697_/X vssd1 vssd1 vccd1 vccd1 _7180_/A sky130_fd_sc_hd__a31o_2
X_8437_ _8437_/A _8437_/B vssd1 vssd1 vccd1 vccd1 _8438_/B sky130_fd_sc_hd__xnor2_1
X_5649_ _6053_/A _6049_/A vssd1 vssd1 vccd1 vccd1 _5695_/B sky130_fd_sc_hd__xnor2_1
X_8368_ _8291_/B _8368_/B vssd1 vssd1 vccd1 vccd1 _8368_/X sky130_fd_sc_hd__and2b_1
XFILLER_104_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7319_ _7297_/A _7048_/B _6728_/A _7293_/A vssd1 vssd1 vccd1 vccd1 _7326_/B sky130_fd_sc_hd__o211a_1
XFILLER_104_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8299_ _8240_/A _8299_/B vssd1 vssd1 vccd1 vccd1 _8299_/X sky130_fd_sc_hd__and2b_1
XFILLER_104_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4951_ _5153_/A _5176_/C _4949_/X _5066_/A vssd1 vssd1 vccd1 vccd1 _4951_/X sky130_fd_sc_hd__o31a_1
X_7670_ _7816_/A _7668_/B _7820_/A vssd1 vssd1 vccd1 vccd1 _7687_/A sky130_fd_sc_hd__a21o_1
XFILLER_51_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4882_ _5235_/A vssd1 vssd1 vccd1 vccd1 _5240_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6621_ _6581_/A _6581_/B _6620_/Y vssd1 vssd1 vccd1 vccd1 _6652_/B sky130_fd_sc_hd__a21o_1
X_6552_ _8699_/Q vssd1 vssd1 vccd1 vccd1 _7511_/S sky130_fd_sc_hd__inv_2
X_6483_ _8700_/Q vssd1 vssd1 vccd1 vccd1 _7514_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5503_ _5486_/A _5486_/B _5502_/Y vssd1 vssd1 vccd1 vccd1 _5507_/B sky130_fd_sc_hd__a21oi_1
X_8222_ _8222_/A _8222_/B vssd1 vssd1 vccd1 vccd1 _8315_/B sky130_fd_sc_hd__xnor2_2
X_5434_ _8650_/Q _5433_/B _5422_/A _5424_/Y vssd1 vssd1 vccd1 vccd1 _5434_/X sky130_fd_sc_hd__a211o_1
X_8153_ _7817_/X _7836_/C _8301_/B vssd1 vssd1 vccd1 vccd1 _8383_/A sky130_fd_sc_hd__o21a_2
XFILLER_87_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7104_ _6728_/A _6905_/B _7048_/X _7060_/A vssd1 vssd1 vccd1 vccd1 _7105_/B sky130_fd_sc_hd__o211ai_2
X_5365_ _5365_/A _5365_/B vssd1 vssd1 vccd1 vccd1 _8639_/D sky130_fd_sc_hd__nor2_1
X_8084_ _8180_/A _8084_/B vssd1 vssd1 vccd1 vccd1 _8086_/B sky130_fd_sc_hd__nand2_1
X_5296_ _5296_/A vssd1 vssd1 vccd1 vccd1 _5296_/X sky130_fd_sc_hd__buf_2
XFILLER_101_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7035_ _7035_/A _7035_/B vssd1 vssd1 vccd1 vccd1 _7036_/B sky130_fd_sc_hd__nor2_1
XFILLER_19_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7937_ _8013_/A _7937_/B vssd1 vssd1 vccd1 vccd1 _7938_/C sky130_fd_sc_hd__nand2_1
XFILLER_35_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7868_ _7867_/B _7867_/C _7867_/A vssd1 vssd1 vccd1 vccd1 _7880_/B sky130_fd_sc_hd__a21o_1
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6819_ _6819_/A _6934_/B vssd1 vssd1 vccd1 vccd1 _6820_/B sky130_fd_sc_hd__xnor2_1
X_7799_ _7902_/A _7933_/B vssd1 vssd1 vccd1 vccd1 _7800_/B sky130_fd_sc_hd__xnor2_1
XFILLER_78_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5150_ _4856_/A _4857_/B _4930_/B vssd1 vssd1 vccd1 vccd1 _5253_/B sky130_fd_sc_hd__a21oi_2
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5081_ _4681_/B _5080_/X _4727_/A vssd1 vssd1 vccd1 vccd1 _5081_/X sky130_fd_sc_hd__o21ba_1
XFILLER_84_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8840_ _8840_/A _4351_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[19] sky130_fd_sc_hd__ebufn_8
X_5983_ _5983_/A _5983_/B vssd1 vssd1 vccd1 vccd1 _5985_/A sky130_fd_sc_hd__nand2_1
XFILLER_25_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7722_ _7722_/A _7722_/B vssd1 vssd1 vccd1 vccd1 _7954_/A sky130_fd_sc_hd__xnor2_1
X_4934_ _4507_/X _5026_/A _4849_/B _5041_/B vssd1 vssd1 vccd1 vccd1 _4955_/B sky130_fd_sc_hd__o31a_1
XFILLER_24_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7653_ _8050_/A vssd1 vssd1 vccd1 vccd1 _8057_/A sky130_fd_sc_hd__clkbuf_2
X_4865_ _4897_/A _4865_/B _4897_/B vssd1 vssd1 vccd1 vccd1 _4990_/B sky130_fd_sc_hd__or3_2
X_6604_ _6592_/A _6584_/B _6561_/B _6556_/X vssd1 vssd1 vccd1 vccd1 _6710_/B sky130_fd_sc_hd__a211o_1
X_7584_ _7627_/A _7583_/X _7541_/X vssd1 vssd1 vccd1 vccd1 _7584_/Y sky130_fd_sc_hd__a21oi_1
X_4796_ _4872_/A _4872_/B _4872_/C vssd1 vssd1 vccd1 vccd1 _4961_/B sky130_fd_sc_hd__nand3_2
XFILLER_21_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6535_ _7545_/B vssd1 vssd1 vccd1 vccd1 _7540_/A sky130_fd_sc_hd__clkbuf_2
X_8205_ _8205_/A _8205_/B _8205_/C vssd1 vssd1 vccd1 vccd1 _8212_/A sky130_fd_sc_hd__and3_1
X_6466_ _8684_/Q _6465_/A _8685_/Q vssd1 vssd1 vccd1 vccd1 _6466_/Y sky130_fd_sc_hd__a21oi_1
X_5417_ _5415_/Y _5417_/B vssd1 vssd1 vccd1 vccd1 _5417_/X sky130_fd_sc_hd__and2b_1
X_6397_ _8670_/Q _8676_/Q _8675_/Q _6397_/D vssd1 vssd1 vccd1 vccd1 _6398_/C sky130_fd_sc_hd__and4bb_1
X_8136_ _8040_/A _8040_/B _8039_/A vssd1 vssd1 vccd1 vccd1 _8194_/B sky130_fd_sc_hd__a21o_1
X_5348_ _5352_/C _5348_/B vssd1 vssd1 vccd1 vccd1 _8634_/D sky130_fd_sc_hd__nor2_1
X_8067_ _8140_/A _8140_/B vssd1 vssd1 vccd1 vccd1 _8071_/A sky130_fd_sc_hd__xnor2_1
XFILLER_101_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7018_ _7018_/A _7018_/B vssd1 vssd1 vccd1 vccd1 _7084_/A sky130_fd_sc_hd__xnor2_2
XFILLER_87_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5279_ _8656_/Q _5271_/X _5278_/X _5273_/X vssd1 vssd1 vccd1 vccd1 _8614_/D sky130_fd_sc_hd__o211a_1
XFILLER_28_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4650_ _4650_/A vssd1 vssd1 vccd1 vccd1 _4784_/A sky130_fd_sc_hd__buf_2
X_6320_ _6320_/A _6326_/A _6326_/B _6326_/C vssd1 vssd1 vccd1 vccd1 _6341_/B sky130_fd_sc_hd__or4_2
X_4581_ _4581_/A _5449_/B vssd1 vssd1 vccd1 vccd1 _4582_/B sky130_fd_sc_hd__nand2_4
X_6251_ _6213_/A _5742_/A _6227_/S _6228_/A _6228_/B vssd1 vssd1 vccd1 vccd1 _6251_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_97_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5202_ _5202_/A _5202_/B _5248_/C _4928_/B vssd1 vssd1 vccd1 vccd1 _5202_/X sky130_fd_sc_hd__or4b_1
X_6182_ _6182_/A _6182_/B vssd1 vssd1 vccd1 vccd1 _6187_/A sky130_fd_sc_hd__nand2_1
XFILLER_96_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5133_ _5175_/B vssd1 vssd1 vccd1 vccd1 _5133_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5064_ _5130_/A vssd1 vssd1 vccd1 vccd1 _5149_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_84_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8823_ _8823_/A _4330_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[2] sky130_fd_sc_hd__ebufn_8
XFILLER_25_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5966_ _6178_/A _6178_/B vssd1 vssd1 vccd1 vccd1 _5967_/B sky130_fd_sc_hd__xor2_1
X_7705_ _7745_/A _7745_/B _7717_/B _7704_/X _7701_/A vssd1 vssd1 vccd1 vccd1 _7740_/B
+ sky130_fd_sc_hd__a311o_4
X_4917_ _5092_/C _4988_/A vssd1 vssd1 vccd1 vccd1 _4946_/A sky130_fd_sc_hd__or2_1
X_8685_ input3/X _8685_/D vssd1 vssd1 vccd1 vccd1 _8685_/Q sky130_fd_sc_hd__dfxtp_1
X_5897_ _5906_/A _5897_/B vssd1 vssd1 vccd1 vccd1 _5898_/B sky130_fd_sc_hd__xnor2_1
X_7636_ _7636_/A _7636_/B vssd1 vssd1 vccd1 vccd1 _7779_/A sky130_fd_sc_hd__xnor2_2
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4848_ _4848_/A _4848_/B vssd1 vssd1 vccd1 vccd1 _5227_/B sky130_fd_sc_hd__nor2_2
XFILLER_32_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7567_ _7593_/B _8707_/Q vssd1 vssd1 vccd1 vccd1 _7594_/A sky130_fd_sc_hd__and2b_1
X_4779_ _4784_/A _4779_/B vssd1 vssd1 vccd1 vccd1 _8610_/D sky130_fd_sc_hd__nor2_1
X_7498_ _7492_/A _7508_/A _7497_/X _7503_/A vssd1 vssd1 vccd1 vccd1 _7498_/Y sky130_fd_sc_hd__o31ai_4
X_6518_ _6514_/A _6511_/X _6513_/X _6517_/X vssd1 vssd1 vccd1 vccd1 _8689_/D sky130_fd_sc_hd__a22o_1
X_6449_ _6450_/B _6450_/C _6448_/Y vssd1 vssd1 vccd1 vccd1 _8678_/D sky130_fd_sc_hd__a21oi_1
X_8119_ _8225_/A _8319_/A _8226_/A vssd1 vssd1 vccd1 vccd1 _8120_/B sky130_fd_sc_hd__o21a_1
XFILLER_57_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5820_ _5820_/A _5820_/B _6218_/A vssd1 vssd1 vccd1 vccd1 _5821_/B sky130_fd_sc_hd__nand3_1
X_5751_ _5849_/B _6185_/A vssd1 vssd1 vccd1 vccd1 _5751_/X sky130_fd_sc_hd__and2_1
X_8470_ _8470_/A _8470_/B vssd1 vssd1 vccd1 vccd1 _8471_/B sky130_fd_sc_hd__xor2_1
X_4702_ _4707_/A _5060_/A vssd1 vssd1 vccd1 vccd1 _4702_/X sky130_fd_sc_hd__or2_1
X_7421_ _7438_/A _7438_/B _7420_/A vssd1 vssd1 vccd1 vccd1 _7424_/A sky130_fd_sc_hd__a21oi_1
X_5682_ _5682_/A _5682_/B vssd1 vssd1 vccd1 vccd1 _5961_/B sky130_fd_sc_hd__or2_2
XFILLER_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4633_ _8586_/Q _4632_/B _4607_/X vssd1 vssd1 vccd1 vccd1 _4634_/B sky130_fd_sc_hd__o21ai_1
X_7352_ _7345_/B _7345_/C _7345_/A vssd1 vssd1 vccd1 vccd1 _7354_/A sky130_fd_sc_hd__o21ba_1
X_4564_ _4564_/A vssd1 vssd1 vccd1 vccd1 _8871_/A sky130_fd_sc_hd__clkbuf_1
X_7283_ _7283_/A _7283_/B vssd1 vssd1 vccd1 vccd1 _7456_/B sky130_fd_sc_hd__xor2_1
X_6303_ _6303_/A _6303_/B _6303_/C vssd1 vssd1 vccd1 vccd1 _6304_/C sky130_fd_sc_hd__nand3_1
XFILLER_89_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4495_ _4495_/A _4495_/B vssd1 vssd1 vccd1 vccd1 _4781_/B sky130_fd_sc_hd__and2_1
X_6234_ _6234_/A _6234_/B vssd1 vssd1 vccd1 vccd1 _6266_/B sky130_fd_sc_hd__xnor2_2
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6165_ _6163_/X _6164_/X _6311_/B vssd1 vssd1 vccd1 vccd1 _6165_/X sky130_fd_sc_hd__o21ba_1
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5116_ _5240_/A _5116_/B _5193_/A _5219_/D vssd1 vssd1 vccd1 vccd1 _5116_/X sky130_fd_sc_hd__or4_1
X_6096_ _6096_/A _6151_/A vssd1 vssd1 vccd1 vccd1 _6099_/A sky130_fd_sc_hd__or2b_1
XFILLER_84_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5047_ _5054_/C _5047_/B _5120_/C _5047_/D vssd1 vssd1 vccd1 vccd1 _5047_/X sky130_fd_sc_hd__or4_1
XFILLER_27_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6998_ _6998_/A _6988_/X vssd1 vssd1 vccd1 vccd1 _7147_/A sky130_fd_sc_hd__or2b_1
XFILLER_80_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5949_ _5949_/A _5949_/B vssd1 vssd1 vccd1 vccd1 _5972_/A sky130_fd_sc_hd__nand2_1
XFILLER_13_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8668_ input3/X _8668_/D vssd1 vssd1 vccd1 vccd1 _8668_/Q sky130_fd_sc_hd__dfxtp_1
X_7619_ _8564_/A _7619_/B vssd1 vssd1 vccd1 vccd1 _7619_/Y sky130_fd_sc_hd__nor2_1
X_8599_ input3/X _8599_/D vssd1 vssd1 vccd1 vccd1 _8599_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7970_ _8023_/B _7969_/C _7969_/A vssd1 vssd1 vccd1 vccd1 _7976_/B sky130_fd_sc_hd__a21o_1
XFILLER_54_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6921_ _6920_/B _7062_/A _6920_/A vssd1 vssd1 vccd1 vccd1 _6922_/C sky130_fd_sc_hd__a21o_1
X_6852_ _6895_/A _6852_/B vssd1 vssd1 vccd1 vccd1 _6854_/B sky130_fd_sc_hd__xnor2_2
XFILLER_81_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5803_ _6214_/A _5803_/B vssd1 vssd1 vccd1 vccd1 _5903_/A sky130_fd_sc_hd__nand2_1
X_6783_ _6954_/B _6881_/A vssd1 vssd1 vccd1 vccd1 _6784_/B sky130_fd_sc_hd__nand2_1
X_8522_ _8522_/A _8522_/B vssd1 vssd1 vccd1 vccd1 _8523_/B sky130_fd_sc_hd__nand2_1
XFILLER_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5734_ _5792_/B _5816_/A vssd1 vssd1 vccd1 vccd1 _5736_/B sky130_fd_sc_hd__xnor2_1
XFILLER_13_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8453_ _8453_/A _8418_/B vssd1 vssd1 vccd1 vccd1 _8453_/X sky130_fd_sc_hd__or2b_1
X_5665_ _5697_/A _5697_/B vssd1 vssd1 vccd1 vccd1 _5746_/A sky130_fd_sc_hd__and2b_1
X_8384_ _8384_/A _8384_/B vssd1 vssd1 vccd1 vccd1 _8445_/B sky130_fd_sc_hd__nand2_1
X_7404_ _7425_/A _7231_/A _7403_/X vssd1 vssd1 vccd1 vccd1 _7422_/B sky130_fd_sc_hd__a21o_1
X_4616_ _4619_/C _4616_/B vssd1 vssd1 vccd1 vccd1 _8580_/D sky130_fd_sc_hd__nor2_1
X_7335_ _7336_/A _7336_/B _7336_/C _7336_/D vssd1 vssd1 vccd1 vccd1 _7337_/B sky130_fd_sc_hd__o22ai_1
X_5596_ _5742_/A _5596_/B vssd1 vssd1 vccd1 vccd1 _5740_/B sky130_fd_sc_hd__xnor2_1
XFILLER_104_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4547_ _4547_/A vssd1 vssd1 vccd1 vccd1 _8867_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_2_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7266_ _7266_/A _7266_/B vssd1 vssd1 vccd1 vccd1 _7270_/A sky130_fd_sc_hd__or2_1
X_4478_ _4478_/A vssd1 vssd1 vccd1 vccd1 _8864_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_104_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7197_ _7223_/A _7197_/B vssd1 vssd1 vccd1 vccd1 _7305_/A sky130_fd_sc_hd__nor2_1
X_6217_ _6217_/A _6217_/B vssd1 vssd1 vccd1 vccd1 _6218_/B sky130_fd_sc_hd__nand2_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6148_ _6300_/A _6300_/B vssd1 vssd1 vccd1 vccd1 _6303_/B sky130_fd_sc_hd__or2_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6079_ _5754_/A _5954_/A _6053_/B _6052_/A vssd1 vssd1 vccd1 vccd1 _6094_/B sky130_fd_sc_hd__a31o_1
XFILLER_18_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8812__90 vssd1 vssd1 vccd1 vccd1 _8812__90/HI _8921_/A sky130_fd_sc_hd__conb_1
XFILLER_72_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5450_ _5449_/B _5449_/C _5615_/A vssd1 vssd1 vccd1 vccd1 _5451_/C sky130_fd_sc_hd__o21ai_1
X_4401_ _4401_/A vssd1 vssd1 vccd1 vccd1 _4401_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5381_ _5462_/B _6346_/A _8661_/Q vssd1 vssd1 vccd1 vccd1 _5381_/X sky130_fd_sc_hd__o21a_1
XFILLER_99_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7120_ _7120_/A _7120_/B vssd1 vssd1 vccd1 vccd1 _7121_/B sky130_fd_sc_hd__xnor2_1
X_4332_ _4333_/A vssd1 vssd1 vccd1 vccd1 _4332_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7051_ _7099_/A _7051_/B _7051_/C vssd1 vssd1 vccd1 vccd1 _7052_/A sky130_fd_sc_hd__or3_1
XFILLER_59_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6002_ _5914_/A _5914_/B _5913_/A vssd1 vssd1 vccd1 vccd1 _6020_/A sky130_fd_sc_hd__a21o_1
XFILLER_82_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7953_ _7889_/A _7865_/B _7865_/C vssd1 vssd1 vccd1 vccd1 _7960_/A sky130_fd_sc_hd__o21bai_1
XFILLER_82_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6904_ _6919_/A _7296_/B _7047_/A vssd1 vssd1 vccd1 vccd1 _6905_/C sky130_fd_sc_hd__and3b_1
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7884_ _7884_/A _7957_/C _7957_/D vssd1 vssd1 vccd1 vccd1 _7972_/A sky130_fd_sc_hd__or3_2
XFILLER_23_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6835_ _8704_/Q _6608_/B vssd1 vssd1 vccd1 vccd1 _6836_/B sky130_fd_sc_hd__or2b_1
XFILLER_62_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6766_ _6766_/A _6829_/B vssd1 vssd1 vccd1 vccd1 _6767_/B sky130_fd_sc_hd__xnor2_1
XFILLER_50_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8505_ _8497_/C _8503_/X _8504_/Y _8501_/B vssd1 vssd1 vccd1 vccd1 _8505_/Y sky130_fd_sc_hd__a2bb2oi_1
X_5717_ _5718_/A _5718_/B vssd1 vssd1 vccd1 vccd1 _5717_/X sky130_fd_sc_hd__or2_1
XFILLER_50_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6697_ _6697_/A _6697_/B _7299_/A vssd1 vssd1 vccd1 vccd1 _6697_/X sky130_fd_sc_hd__and3_1
XFILLER_40_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8436_ _8421_/A _8421_/B _8435_/Y vssd1 vssd1 vccd1 vccd1 _8438_/A sky130_fd_sc_hd__a21bo_1
X_5648_ _5671_/A _5980_/A vssd1 vssd1 vccd1 vccd1 _6049_/A sky130_fd_sc_hd__nor2_1
XFILLER_40_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8367_ _8442_/A _8442_/B vssd1 vssd1 vccd1 vccd1 _8370_/A sky130_fd_sc_hd__xnor2_1
X_5579_ _5595_/B vssd1 vssd1 vccd1 vccd1 _5731_/A sky130_fd_sc_hd__clkbuf_2
X_8298_ _8298_/A _8298_/B vssd1 vssd1 vccd1 vccd1 _8347_/A sky130_fd_sc_hd__xor2_1
X_7318_ _7318_/A _7318_/B vssd1 vssd1 vccd1 vccd1 _7326_/A sky130_fd_sc_hd__xnor2_2
X_7249_ _7293_/A _7249_/B _7294_/A vssd1 vssd1 vccd1 vccd1 _7317_/B sky130_fd_sc_hd__and3_1
XFILLER_49_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8789__67 vssd1 vssd1 vccd1 vccd1 _8789__67/HI _8898_/A sky130_fd_sc_hd__conb_1
XFILLER_58_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4950_ _5231_/A vssd1 vssd1 vccd1 vccd1 _5066_/A sky130_fd_sc_hd__clkbuf_2
X_4881_ _5153_/A _5199_/A vssd1 vssd1 vccd1 vccd1 _4881_/X sky130_fd_sc_hd__or2_1
X_6620_ _6620_/A _6660_/B vssd1 vssd1 vccd1 vccd1 _6620_/Y sky130_fd_sc_hd__nand2_1
XFILLER_32_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6551_ _8595_/Q _8699_/Q vssd1 vssd1 vccd1 vccd1 _6592_/A sky130_fd_sc_hd__nand2b_4
X_5502_ _8662_/Q _7688_/B _5482_/B vssd1 vssd1 vccd1 vccd1 _5502_/Y sky130_fd_sc_hd__o21ai_1
X_6482_ _8701_/Q vssd1 vssd1 vccd1 vccd1 _7518_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_8221_ _8229_/A _8406_/B vssd1 vssd1 vccd1 vccd1 _8222_/B sky130_fd_sc_hd__xor2_1
X_5433_ _8651_/Q _5433_/B vssd1 vssd1 vccd1 vccd1 _5437_/B sky130_fd_sc_hd__or2_1
X_8152_ _8152_/A vssd1 vssd1 vccd1 vccd1 _8301_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5364_ _8639_/Q _5366_/C _5357_/X vssd1 vssd1 vccd1 vccd1 _5365_/B sky130_fd_sc_hd__o21ai_1
X_7103_ _7103_/A _7103_/B vssd1 vssd1 vccd1 vccd1 _7105_/A sky130_fd_sc_hd__nand2_1
XFILLER_101_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8083_ _8083_/A _8083_/B vssd1 vssd1 vccd1 vccd1 _8084_/B sky130_fd_sc_hd__or2_1
X_5295_ _8621_/Q _5300_/B vssd1 vssd1 vccd1 vccd1 _5295_/X sky130_fd_sc_hd__or2_1
XFILLER_101_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7034_ _7034_/A _7034_/B vssd1 vssd1 vccd1 vccd1 _7035_/B sky130_fd_sc_hd__nor2_1
XFILLER_19_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7936_ _7936_/A _7936_/B vssd1 vssd1 vccd1 vccd1 _7937_/B sky130_fd_sc_hd__nand2_1
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7867_ _7867_/A _7867_/B _7867_/C vssd1 vssd1 vccd1 vccd1 _7880_/A sky130_fd_sc_hd__nand3_1
XFILLER_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6818_ _6899_/A _7023_/A vssd1 vssd1 vccd1 vccd1 _6934_/B sky130_fd_sc_hd__xor2_1
X_7798_ _7904_/C _7798_/B vssd1 vssd1 vccd1 vccd1 _7933_/B sky130_fd_sc_hd__xor2_1
XFILLER_50_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6749_ _6719_/A _6700_/B _6769_/A vssd1 vssd1 vccd1 vccd1 _6768_/B sky130_fd_sc_hd__a21bo_1
X_8419_ _8419_/A _8419_/B vssd1 vssd1 vccd1 vccd1 _8435_/B sky130_fd_sc_hd__xnor2_1
XFILLER_2_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5080_ _5243_/A _5074_/X _5075_/Y _4789_/A _5079_/X vssd1 vssd1 vccd1 vccd1 _5080_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_2_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5982_ _6183_/A _5982_/B vssd1 vssd1 vccd1 vccd1 _5988_/A sky130_fd_sc_hd__xnor2_2
X_7721_ _7887_/A _8118_/A vssd1 vssd1 vccd1 vccd1 _7777_/C sky130_fd_sc_hd__or2_1
X_4933_ _4933_/A vssd1 vssd1 vccd1 vccd1 _5231_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7652_ _7796_/A vssd1 vssd1 vccd1 vccd1 _8050_/A sky130_fd_sc_hd__buf_2
X_4864_ _5227_/B _4864_/B vssd1 vssd1 vccd1 vccd1 _4866_/A sky130_fd_sc_hd__nand2_1
XFILLER_20_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6603_ _6605_/B _8702_/Q vssd1 vssd1 vccd1 vccd1 _6712_/A sky130_fd_sc_hd__or2b_1
X_7583_ _8568_/A vssd1 vssd1 vccd1 vccd1 _7583_/X sky130_fd_sc_hd__clkbuf_2
X_4795_ _5620_/A _4795_/B vssd1 vssd1 vccd1 vccd1 _4872_/C sky130_fd_sc_hd__xnor2_2
X_6534_ _6533_/A _6540_/A _6533_/C vssd1 vssd1 vccd1 vccd1 _6534_/X sky130_fd_sc_hd__a21o_1
X_6465_ _6465_/A _6465_/B vssd1 vssd1 vccd1 vccd1 _8683_/D sky130_fd_sc_hd__nor2_1
X_8204_ _8138_/A _8138_/B _8203_/X vssd1 vssd1 vccd1 vccd1 _8240_/A sky130_fd_sc_hd__a21oi_2
X_5416_ _5607_/A _5416_/B vssd1 vssd1 vccd1 vccd1 _5417_/B sky130_fd_sc_hd__nand2_1
X_6396_ _8674_/Q _8678_/Q _8677_/Q _8673_/Q vssd1 vssd1 vccd1 vccd1 _6398_/B sky130_fd_sc_hd__and4bb_1
X_8135_ _8031_/A _8317_/B _8462_/B vssd1 vssd1 vccd1 vccd1 _8398_/A sky130_fd_sc_hd__a21o_2
X_5347_ _8634_/Q _5346_/B _5325_/X vssd1 vssd1 vccd1 vccd1 _5348_/B sky130_fd_sc_hd__o21ai_1
XFILLER_101_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8066_ _8066_/A _8066_/B vssd1 vssd1 vccd1 vccd1 _8140_/B sky130_fd_sc_hd__nor2_1
X_5278_ _8614_/Q _5288_/B vssd1 vssd1 vccd1 vccd1 _5278_/X sky130_fd_sc_hd__or2_1
X_7017_ _7142_/B _7017_/B vssd1 vssd1 vccd1 vccd1 _7018_/B sky130_fd_sc_hd__xnor2_1
XFILLER_46_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8759__37 vssd1 vssd1 vccd1 vccd1 _8759__37/HI _8854_/A sky130_fd_sc_hd__conb_1
XFILLER_83_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7919_ _7920_/A _7920_/B vssd1 vssd1 vccd1 vccd1 _8006_/B sky130_fd_sc_hd__nor2_1
XFILLER_43_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8899_ _8899_/A _4413_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[8] sky130_fd_sc_hd__ebufn_8
XFILLER_51_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8773__51 vssd1 vssd1 vccd1 vccd1 _8773__51/HI _8882_/A sky130_fd_sc_hd__conb_1
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4580_ _8591_/Q _5406_/B vssd1 vssd1 vccd1 vccd1 _5449_/B sky130_fd_sc_hd__nand2_2
X_6250_ _6222_/A _6222_/B _6249_/Y vssd1 vssd1 vccd1 vccd1 _6262_/A sky130_fd_sc_hd__o21a_1
XFILLER_103_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6181_ _5754_/B _6204_/A _5988_/B _5988_/A vssd1 vssd1 vccd1 vccd1 _6188_/A sky130_fd_sc_hd__a22oi_2
X_5201_ _5054_/D _5047_/D _5044_/D vssd1 vssd1 vccd1 vccd1 _5201_/X sky130_fd_sc_hd__o21a_1
XFILLER_69_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5132_ _5243_/A _5132_/B _5159_/C vssd1 vssd1 vccd1 vccd1 _5132_/X sky130_fd_sc_hd__or3_1
XFILLER_96_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5063_ _5172_/A _5135_/D vssd1 vssd1 vccd1 vccd1 _5130_/A sky130_fd_sc_hd__or2_1
XFILLER_37_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8822_ _8822_/A _4329_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[1] sky130_fd_sc_hd__ebufn_8
XFILLER_37_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5965_ _5956_/B _5965_/B _6182_/B vssd1 vssd1 vccd1 vccd1 _6178_/B sky130_fd_sc_hd__and3b_1
XFILLER_25_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7704_ _7702_/Y _6605_/B _6560_/B _8538_/A vssd1 vssd1 vccd1 vccd1 _7704_/X sky130_fd_sc_hd__o211a_1
XFILLER_52_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4916_ _5159_/B _4916_/B vssd1 vssd1 vccd1 vccd1 _4988_/A sky130_fd_sc_hd__or2_1
X_8684_ input3/X _8684_/D vssd1 vssd1 vccd1 vccd1 _8684_/Q sky130_fd_sc_hd__dfxtp_1
X_5896_ _5896_/A _5896_/B vssd1 vssd1 vccd1 vccd1 _5900_/B sky130_fd_sc_hd__and2_1
X_7635_ _7633_/X _7643_/A vssd1 vssd1 vccd1 vccd1 _7636_/B sky130_fd_sc_hd__and2b_1
X_4847_ _4847_/A vssd1 vssd1 vccd1 vccd1 _5041_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7566_ _8710_/Q vssd1 vssd1 vccd1 vccd1 _7593_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_20_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4778_ _4781_/A _4778_/B vssd1 vssd1 vccd1 vccd1 _4779_/B sky130_fd_sc_hd__xor2_1
X_7497_ _7494_/Y _7505_/C _7492_/D _7492_/C _7474_/X vssd1 vssd1 vccd1 vccd1 _7497_/X
+ sky130_fd_sc_hd__a2111o_1
X_6517_ _6515_/Y _6517_/B vssd1 vssd1 vccd1 vccd1 _6517_/X sky130_fd_sc_hd__and2b_1
X_6448_ _6450_/B _6450_/C _6409_/B vssd1 vssd1 vccd1 vccd1 _6448_/Y sky130_fd_sc_hd__o21ai_1
X_6379_ _6379_/A _6379_/B vssd1 vssd1 vccd1 vccd1 _8664_/D sky130_fd_sc_hd__nor2_1
X_8118_ _8118_/A _8317_/B vssd1 vssd1 vccd1 vccd1 _8226_/A sky130_fd_sc_hd__or2_1
XFILLER_88_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8049_ _8301_/A _8060_/B vssd1 vssd1 vccd1 vccd1 _8280_/A sky130_fd_sc_hd__nand2_1
XFILLER_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5750_ _5953_/B _5957_/B vssd1 vssd1 vccd1 vccd1 _6185_/A sky130_fd_sc_hd__or2_2
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5681_ _5680_/A _5680_/B _5680_/C vssd1 vssd1 vccd1 vccd1 _5682_/B sky130_fd_sc_hd__a21oi_1
X_4701_ _4701_/A vssd1 vssd1 vccd1 vccd1 _5060_/A sky130_fd_sc_hd__clkbuf_2
X_7420_ _7420_/A _7420_/B vssd1 vssd1 vccd1 vccd1 _7438_/B sky130_fd_sc_hd__nor2_1
X_4632_ _8586_/Q _4632_/B vssd1 vssd1 vccd1 vccd1 _4637_/C sky130_fd_sc_hd__and2_1
XFILLER_30_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7351_ _7343_/A _7343_/B _7350_/X vssd1 vssd1 vccd1 vccd1 _7355_/A sky130_fd_sc_hd__o21a_1
X_4563_ _8617_/Q _4563_/B vssd1 vssd1 vccd1 vccd1 _4564_/A sky130_fd_sc_hd__and2_1
X_7282_ _7282_/A _7282_/B vssd1 vssd1 vccd1 vccd1 _7283_/B sky130_fd_sc_hd__xnor2_1
X_4494_ _4775_/A _4769_/A _4535_/C vssd1 vssd1 vccd1 vccd1 _4495_/B sky130_fd_sc_hd__and3_1
X_6302_ _6302_/A _6302_/B vssd1 vssd1 vccd1 vccd1 _6337_/A sky130_fd_sc_hd__xnor2_1
XFILLER_89_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6233_ _6233_/A _6233_/B vssd1 vssd1 vccd1 vccd1 _6234_/B sky130_fd_sc_hd__xor2_2
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6164_ _6303_/A _6163_/A _6164_/C _6164_/D vssd1 vssd1 vccd1 vccd1 _6164_/X sky130_fd_sc_hd__and4bb_1
XFILLER_97_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5115_ _5119_/B _5115_/B vssd1 vssd1 vccd1 vccd1 _5115_/X sky130_fd_sc_hd__or2_1
X_6095_ _6096_/A _6095_/B _6095_/C vssd1 vssd1 vccd1 vccd1 _6151_/A sky130_fd_sc_hd__or3_1
XFILLER_69_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5046_ _5046_/A _5046_/B vssd1 vssd1 vccd1 vccd1 _5047_/D sky130_fd_sc_hd__or2_1
XFILLER_27_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6997_ _6987_/A _6987_/B _6996_/X vssd1 vssd1 vccd1 vccd1 _7086_/A sky130_fd_sc_hd__a21oi_2
XFILLER_53_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5948_ _5875_/A _5875_/B _5876_/B _5920_/B vssd1 vssd1 vccd1 vccd1 _5975_/A sky130_fd_sc_hd__o22a_1
XFILLER_25_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8667_ input3/X _8667_/D vssd1 vssd1 vccd1 vccd1 _8667_/Q sky130_fd_sc_hd__dfxtp_1
X_5879_ _5879_/A _5896_/A _5879_/C vssd1 vssd1 vccd1 vccd1 _5887_/A sky130_fd_sc_hd__and3_1
X_7618_ _7618_/A _7618_/B vssd1 vssd1 vccd1 vccd1 _7619_/B sky130_fd_sc_hd__xnor2_1
X_8598_ input3/X _8598_/D vssd1 vssd1 vccd1 vccd1 _8598_/Q sky130_fd_sc_hd__dfxtp_1
X_7549_ _8724_/Q vssd1 vssd1 vccd1 vccd1 _8561_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_5_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8743__21 vssd1 vssd1 vccd1 vccd1 _8743__21/HI _8838_/A sky130_fd_sc_hd__conb_1
XFILLER_31_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6920_ _6920_/A _6920_/B _7062_/A vssd1 vssd1 vccd1 vccd1 _7062_/B sky130_fd_sc_hd__nand3_1
X_6851_ _6851_/A _6851_/B vssd1 vssd1 vccd1 vccd1 _6852_/B sky130_fd_sc_hd__xor2_2
XFILLER_62_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5802_ _6215_/A _5800_/X _5907_/A _5803_/B vssd1 vssd1 vccd1 vccd1 _6220_/B sky130_fd_sc_hd__o22a_2
X_6782_ _6954_/B _6881_/A vssd1 vssd1 vccd1 vccd1 _6886_/A sky130_fd_sc_hd__or2_1
X_8521_ _8522_/A _8522_/B vssd1 vssd1 vccd1 vccd1 _8526_/S sky130_fd_sc_hd__or2_1
XFILLER_62_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5733_ _5589_/A _5589_/B _5587_/Y vssd1 vssd1 vccd1 vccd1 _5816_/A sky130_fd_sc_hd__a21oi_1
X_8452_ _8418_/B _8453_/A vssd1 vssd1 vccd1 vccd1 _8452_/X sky130_fd_sc_hd__and2b_1
X_5664_ _5704_/A _5706_/A vssd1 vssd1 vccd1 vccd1 _5697_/B sky130_fd_sc_hd__xnor2_1
X_8383_ _8383_/A _8384_/B _8445_/C vssd1 vssd1 vccd1 vccd1 _8472_/A sky130_fd_sc_hd__and3_1
X_7403_ _7236_/A _6876_/A _7137_/X vssd1 vssd1 vccd1 vccd1 _7403_/X sky130_fd_sc_hd__o21a_1
X_4615_ _8580_/Q _4614_/B _4595_/X vssd1 vssd1 vccd1 vccd1 _4616_/B sky130_fd_sc_hd__o21ai_1
X_5595_ _5595_/A _5595_/B vssd1 vssd1 vccd1 vccd1 _5596_/B sky130_fd_sc_hd__xor2_1
X_7334_ _7270_/A _7313_/B _7334_/C _7334_/D vssd1 vssd1 vccd1 vccd1 _7336_/A sky130_fd_sc_hd__and4bb_1
X_4546_ _8613_/Q _4552_/B vssd1 vssd1 vccd1 vccd1 _4547_/A sky130_fd_sc_hd__and2_1
XFILLER_104_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7265_ _7265_/A _7265_/B vssd1 vssd1 vccd1 vccd1 _7266_/B sky130_fd_sc_hd__and2_1
X_4477_ _4520_/A _4709_/A vssd1 vssd1 vccd1 vccd1 _4478_/A sky130_fd_sc_hd__or2_1
XFILLER_89_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7196_ _7223_/B _7289_/B vssd1 vssd1 vccd1 vccd1 _7196_/X sky130_fd_sc_hd__and2b_1
X_6216_ _6215_/B _6215_/C _6215_/A vssd1 vssd1 vccd1 vccd1 _6217_/B sky130_fd_sc_hd__a21oi_1
X_6147_ _6302_/A _6302_/B vssd1 vssd1 vccd1 vccd1 _6300_/B sky130_fd_sc_hd__or2b_1
XFILLER_38_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6078_ _6046_/Y _6108_/A _6054_/B vssd1 vssd1 vccd1 vccd1 _6087_/B sky130_fd_sc_hd__a21bo_1
X_5029_ _5083_/A _5029_/B _5241_/C _5215_/C vssd1 vssd1 vccd1 vccd1 _5029_/X sky130_fd_sc_hd__or4_1
XFILLER_26_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8719_ input3/X _8719_/D vssd1 vssd1 vccd1 vccd1 _8719_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4400_ _4401_/A vssd1 vssd1 vccd1 vccd1 _4400_/Y sky130_fd_sc_hd__inv_2
X_5380_ _8659_/Q vssd1 vssd1 vccd1 vccd1 _6346_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4331_ _4333_/A vssd1 vssd1 vccd1 vccd1 _4331_/Y sky130_fd_sc_hd__inv_2
X_7050_ _7060_/A _7060_/C _7049_/Y vssd1 vssd1 vccd1 vccd1 _7051_/C sky130_fd_sc_hd__a21oi_1
XFILLER_101_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6001_ _6001_/A _6207_/B vssd1 vssd1 vccd1 vccd1 _6021_/A sky130_fd_sc_hd__and2_1
XFILLER_94_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7952_ _7880_/B _7880_/C _7880_/A vssd1 vssd1 vccd1 vccd1 _7969_/A sky130_fd_sc_hd__a21bo_1
X_6903_ _6919_/A _7245_/B _7048_/C _6798_/B vssd1 vssd1 vccd1 vccd1 _6905_/B sky130_fd_sc_hd__o22a_1
X_7883_ _7882_/B _7882_/C _7882_/A vssd1 vssd1 vccd1 vccd1 _7894_/B sky130_fd_sc_hd__a21o_1
XFILLER_35_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6834_ _6834_/A _6834_/B vssd1 vssd1 vccd1 vccd1 _6942_/A sky130_fd_sc_hd__xnor2_1
X_6765_ _7020_/A _6765_/B vssd1 vssd1 vccd1 vccd1 _6829_/B sky130_fd_sc_hd__xnor2_1
XFILLER_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8504_ _8500_/B _8500_/C _8500_/A vssd1 vssd1 vccd1 vccd1 _8504_/Y sky130_fd_sc_hd__o21ai_1
X_5716_ _5603_/A _5603_/B _5715_/X vssd1 vssd1 vccd1 vccd1 _5745_/A sky130_fd_sc_hd__a21oi_2
XFILLER_31_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8435_ _8435_/A _8435_/B vssd1 vssd1 vccd1 vccd1 _8435_/Y sky130_fd_sc_hd__nand2_1
X_6696_ _7418_/B _6697_/B _7293_/B _6697_/A vssd1 vssd1 vccd1 vccd1 _7167_/B sky130_fd_sc_hd__a22o_1
XFILLER_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5647_ _5647_/A _5647_/B vssd1 vssd1 vccd1 vccd1 _5980_/A sky130_fd_sc_hd__xor2_2
X_8366_ _8441_/A _8366_/B vssd1 vssd1 vccd1 vccd1 _8442_/B sky130_fd_sc_hd__xnor2_1
X_5578_ _5578_/A _5578_/B vssd1 vssd1 vccd1 vccd1 _5721_/A sky130_fd_sc_hd__nand2_1
X_8297_ _8297_/A _8353_/B vssd1 vssd1 vccd1 vccd1 _8298_/B sky130_fd_sc_hd__xnor2_1
X_7317_ _7317_/A _7317_/B vssd1 vssd1 vccd1 vccd1 _7318_/A sky130_fd_sc_hd__xnor2_1
X_4529_ _8593_/Q _5083_/A vssd1 vssd1 vccd1 vccd1 _5214_/A sky130_fd_sc_hd__or2_1
XFILLER_104_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7248_ _7296_/C _7248_/B vssd1 vssd1 vccd1 vccd1 _7317_/A sky130_fd_sc_hd__xor2_1
X_7179_ _7179_/A _7239_/B vssd1 vssd1 vccd1 vccd1 _7182_/A sky130_fd_sc_hd__or2b_1
XFILLER_85_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4880_ _5130_/B vssd1 vssd1 vccd1 vccd1 _5199_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_44_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6550_ _6550_/A vssd1 vssd1 vccd1 vccd1 _8694_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5501_ _6608_/B _6371_/A vssd1 vssd1 vccd1 vccd1 _5507_/A sky130_fd_sc_hd__and2b_1
X_6481_ _7545_/A _6505_/A _7537_/B vssd1 vssd1 vccd1 vccd1 _6481_/Y sky130_fd_sc_hd__o21ai_1
X_8220_ _7757_/B _8331_/B _8113_/B _8205_/B vssd1 vssd1 vccd1 vccd1 _8315_/A sky130_fd_sc_hd__a22o_1
X_5432_ _5447_/A _5433_/B vssd1 vssd1 vccd1 vccd1 _5442_/A sky130_fd_sc_hd__nand2_1
XFILLER_99_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8151_ _8151_/A _8151_/B vssd1 vssd1 vccd1 vccd1 _8155_/A sky130_fd_sc_hd__xor2_1
X_5363_ _8639_/Q _5366_/C vssd1 vssd1 vccd1 vccd1 _5365_/A sky130_fd_sc_hd__and2_1
X_7102_ _7115_/B _7101_/B _7101_/C _7101_/D vssd1 vssd1 vccd1 vccd1 _7103_/B sky130_fd_sc_hd__a22o_1
X_8082_ _8083_/A _8083_/B vssd1 vssd1 vccd1 vccd1 _8180_/A sky130_fd_sc_hd__nand2_1
X_5294_ _8695_/Q _5285_/X _5293_/X _5283_/X vssd1 vssd1 vccd1 vccd1 _8620_/D sky130_fd_sc_hd__o211a_1
XFILLER_101_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7033_ _7034_/A _7034_/B vssd1 vssd1 vccd1 vccd1 _7035_/A sky130_fd_sc_hd__and2_1
XFILLER_101_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7935_ _7936_/A _7936_/B vssd1 vssd1 vccd1 vccd1 _8013_/A sky130_fd_sc_hd__or2_1
XFILLER_35_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7866_ _7865_/B _7865_/C _7889_/A vssd1 vssd1 vccd1 vccd1 _7867_/C sky130_fd_sc_hd__o21ai_1
XFILLER_23_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6817_ _6949_/A vssd1 vssd1 vccd1 vccd1 _7023_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7797_ _7682_/A _7995_/B _7796_/X vssd1 vssd1 vccd1 vccd1 _7798_/B sky130_fd_sc_hd__o21a_1
XFILLER_50_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6748_ _6868_/A _6748_/B vssd1 vssd1 vccd1 vccd1 _7185_/A sky130_fd_sc_hd__and2_1
XFILLER_51_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6679_ _7237_/C vssd1 vssd1 vccd1 vccd1 _7048_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_8418_ _8453_/A _8418_/B vssd1 vssd1 vccd1 vccd1 _8419_/B sky130_fd_sc_hd__xnor2_1
X_8349_ _8349_/A _8352_/B vssd1 vssd1 vccd1 vccd1 _8429_/B sky130_fd_sc_hd__xnor2_1
XFILLER_2_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5981_ _5754_/A _5986_/A _5980_/X vssd1 vssd1 vccd1 vccd1 _5982_/B sky130_fd_sc_hd__o21a_1
X_7720_ _8116_/C vssd1 vssd1 vccd1 vccd1 _8118_/A sky130_fd_sc_hd__clkbuf_2
X_4932_ _4990_/A _5175_/B vssd1 vssd1 vccd1 vccd1 _4941_/C sky130_fd_sc_hd__nand2_1
X_7651_ _7666_/A _7790_/A vssd1 vssd1 vccd1 vccd1 _7651_/Y sky130_fd_sc_hd__nand2_1
X_6602_ _7529_/A _7688_/B vssd1 vssd1 vccd1 vccd1 _6837_/A sky130_fd_sc_hd__nand2_1
X_4863_ _5119_/B _5072_/B vssd1 vssd1 vccd1 vccd1 _5241_/B sky130_fd_sc_hd__or2_1
XFILLER_20_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7582_ _8535_/S vssd1 vssd1 vccd1 vccd1 _8568_/A sky130_fd_sc_hd__clkbuf_2
X_4794_ _4848_/B _4794_/B vssd1 vssd1 vccd1 vccd1 _4872_/B sky130_fd_sc_hd__nand2_1
XFILLER_20_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6533_ _6533_/A _6540_/A _6533_/C vssd1 vssd1 vccd1 vccd1 _6545_/A sky130_fd_sc_hd__nand3_1
XFILLER_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6464_ _8683_/Q _6463_/B _6419_/X vssd1 vssd1 vccd1 vccd1 _6465_/B sky130_fd_sc_hd__o21ai_1
X_8203_ _8133_/A _8203_/B vssd1 vssd1 vccd1 vccd1 _8203_/X sky130_fd_sc_hd__and2b_1
X_5415_ _5607_/A _5416_/B vssd1 vssd1 vccd1 vccd1 _5415_/Y sky130_fd_sc_hd__nor2_1
X_6395_ _8668_/Q _8672_/Q _6430_/A _8667_/Q vssd1 vssd1 vccd1 vccd1 _6400_/B sky130_fd_sc_hd__and4bb_1
X_8134_ _8134_/A _8134_/B vssd1 vssd1 vccd1 vccd1 _8462_/B sky130_fd_sc_hd__nor2_2
X_5346_ _8634_/Q _5346_/B vssd1 vssd1 vccd1 vccd1 _5352_/C sky130_fd_sc_hd__and2_1
XFILLER_87_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8065_ _8065_/A _8437_/A vssd1 vssd1 vccd1 vccd1 _8066_/B sky130_fd_sc_hd__xnor2_1
X_5277_ _5290_/A vssd1 vssd1 vccd1 vccd1 _5288_/B sky130_fd_sc_hd__clkbuf_2
X_7016_ _7202_/A _7016_/B vssd1 vssd1 vccd1 vccd1 _7017_/B sky130_fd_sc_hd__xnor2_2
XFILLER_87_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7918_ _7904_/C _7798_/B _7682_/A _7995_/B vssd1 vssd1 vccd1 vccd1 _7920_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_70_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8898_ _8898_/A _4411_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[7] sky130_fd_sc_hd__ebufn_8
X_7849_ _7849_/A _7849_/B vssd1 vssd1 vccd1 vccd1 _8522_/A sky130_fd_sc_hd__nand2_1
XFILLER_23_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6180_ _6180_/A _6180_/B vssd1 vssd1 vccd1 vccd1 _6204_/A sky130_fd_sc_hd__nor2_1
X_5200_ _5075_/Y _5193_/Y _5192_/Y _5144_/B _5057_/A vssd1 vssd1 vccd1 vccd1 _5200_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5131_ _5137_/C vssd1 vssd1 vccd1 vccd1 _5159_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_69_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5062_ _5214_/B _5214_/C _5240_/C _5239_/B vssd1 vssd1 vccd1 vccd1 _5062_/X sky130_fd_sc_hd__or4_1
XFILLER_96_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8821_ _8821_/A _4459_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[0] sky130_fd_sc_hd__ebufn_8
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7703_ _8539_/A vssd1 vssd1 vccd1 vccd1 _8538_/A sky130_fd_sc_hd__inv_2
X_5964_ _5753_/A _5964_/B _6182_/A vssd1 vssd1 vccd1 vccd1 _6182_/B sky130_fd_sc_hd__nand3b_1
X_4915_ _4989_/A vssd1 vssd1 vccd1 vccd1 _5071_/A sky130_fd_sc_hd__clkbuf_2
X_8683_ input3/X _8683_/D vssd1 vssd1 vccd1 vccd1 _8683_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5895_ _5895_/A _5895_/B vssd1 vssd1 vccd1 vccd1 _5900_/A sky130_fd_sc_hd__and2_1
X_7634_ _7634_/A _7593_/B vssd1 vssd1 vccd1 vccd1 _7643_/A sky130_fd_sc_hd__or2b_2
X_4846_ _4849_/A _4850_/B _4909_/A _4850_/A vssd1 vssd1 vccd1 vccd1 _4847_/A sky130_fd_sc_hd__or4b_1
X_7565_ _8713_/Q vssd1 vssd1 vccd1 vccd1 _7616_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6516_ _6567_/A _6516_/B vssd1 vssd1 vccd1 vccd1 _6517_/B sky130_fd_sc_hd__nand2_1
X_4777_ _4777_/A vssd1 vssd1 vccd1 vccd1 _8609_/D sky130_fd_sc_hd__clkbuf_1
X_7496_ _7496_/A _7496_/B vssd1 vssd1 vccd1 vccd1 _7505_/C sky130_fd_sc_hd__nor2_1
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6447_ _6450_/C _6447_/B vssd1 vssd1 vccd1 vccd1 _8677_/D sky130_fd_sc_hd__nor2_1
X_6378_ _8664_/Q _5419_/A _6376_/X _4650_/A vssd1 vssd1 vccd1 vccd1 _6379_/B sky130_fd_sc_hd__a31o_1
XFILLER_102_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8819__97 vssd1 vssd1 vccd1 vccd1 _8819__97/HI _8928_/A sky130_fd_sc_hd__conb_1
X_8117_ _8395_/B _8230_/A _8117_/S vssd1 vssd1 vccd1 vccd1 _8319_/A sky130_fd_sc_hd__mux2_1
X_5329_ _6475_/B _5330_/C _5328_/Y vssd1 vssd1 vccd1 vccd1 _8628_/D sky130_fd_sc_hd__a21oi_1
X_8048_ _8103_/A _8103_/B vssd1 vssd1 vccd1 vccd1 _8072_/A sky130_fd_sc_hd__xor2_1
XFILLER_16_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5680_ _5680_/A _5680_/B _5680_/C vssd1 vssd1 vccd1 vccd1 _5682_/A sky130_fd_sc_hd__and3_1
X_4700_ _4994_/A _4994_/B vssd1 vssd1 vccd1 vccd1 _4701_/A sky130_fd_sc_hd__nor2_1
XFILLER_8_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4631_ _4631_/A vssd1 vssd1 vccd1 vccd1 _8585_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7350_ _7350_/A _7350_/B vssd1 vssd1 vccd1 vccd1 _7350_/X sky130_fd_sc_hd__or2_1
X_4562_ _4562_/A vssd1 vssd1 vccd1 vccd1 _8870_/A sky130_fd_sc_hd__clkbuf_1
X_7281_ _7362_/A _7362_/B _7280_/X vssd1 vssd1 vccd1 vccd1 _7283_/A sky130_fd_sc_hd__a21o_1
X_4493_ _5620_/A vssd1 vssd1 vccd1 vccd1 _4535_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_6301_ _6303_/B _6301_/B vssd1 vssd1 vccd1 vccd1 _6301_/X sky130_fd_sc_hd__and2_1
XFILLER_103_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6232_ _6232_/A _6232_/B vssd1 vssd1 vccd1 vccd1 _6233_/B sky130_fd_sc_hd__nor2_1
XFILLER_69_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6163_ _6163_/A _6164_/D vssd1 vssd1 vccd1 vccd1 _6163_/X sky130_fd_sc_hd__and2_1
XFILLER_85_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5114_ _5194_/A _5114_/B vssd1 vssd1 vccd1 vccd1 _5248_/C sky130_fd_sc_hd__nand2_1
X_6094_ _6094_/A _6094_/B vssd1 vssd1 vccd1 vccd1 _6095_/C sky130_fd_sc_hd__xor2_1
XFILLER_97_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5045_ _5045_/A _5166_/B vssd1 vssd1 vccd1 vccd1 _5120_/C sky130_fd_sc_hd__or2_1
XFILLER_84_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6996_ _6986_/B _6996_/B vssd1 vssd1 vccd1 vccd1 _6996_/X sky130_fd_sc_hd__and2b_1
X_5947_ _5939_/A _5939_/B _5946_/Y vssd1 vssd1 vccd1 vccd1 _6171_/B sky130_fd_sc_hd__a21o_1
XFILLER_40_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8666_ input3/X _8666_/D vssd1 vssd1 vccd1 vccd1 _8666_/Q sky130_fd_sc_hd__dfxtp_1
X_7617_ _7617_/A _7621_/B vssd1 vssd1 vccd1 vccd1 _7618_/B sky130_fd_sc_hd__nand2_1
X_5878_ _5822_/A _5822_/B _5877_/X vssd1 vssd1 vccd1 vccd1 _5917_/A sky130_fd_sc_hd__a21oi_2
X_4829_ _4829_/A _4857_/B vssd1 vssd1 vccd1 vccd1 _4829_/Y sky130_fd_sc_hd__nor2_1
XFILLER_21_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8597_ input3/X _8597_/D vssd1 vssd1 vccd1 vccd1 _8597_/Q sky130_fd_sc_hd__dfxtp_2
X_7548_ _7548_/A vssd1 vssd1 vccd1 vccd1 _8705_/D sky130_fd_sc_hd__clkbuf_1
X_7479_ _7479_/A _7479_/B vssd1 vssd1 vccd1 vccd1 _7486_/A sky130_fd_sc_hd__xnor2_1
XFILLER_4_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6850_ _6850_/A _6970_/B vssd1 vssd1 vccd1 vccd1 _6851_/B sky130_fd_sc_hd__xnor2_2
XFILLER_81_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6781_ _6863_/A _6869_/A vssd1 vssd1 vccd1 vccd1 _6881_/A sky130_fd_sc_hd__or2_1
XFILLER_62_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5801_ _5883_/A _6034_/B _5801_/C vssd1 vssd1 vccd1 vccd1 _5907_/A sky130_fd_sc_hd__and3b_1
X_8520_ _8520_/A _8520_/B vssd1 vssd1 vccd1 vccd1 _8522_/B sky130_fd_sc_hd__nor2_1
XFILLER_50_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5732_ _5595_/A _5803_/B _5596_/B _5895_/A vssd1 vssd1 vccd1 vccd1 _5736_/A sky130_fd_sc_hd__a22o_1
X_8451_ _8451_/A _8451_/B vssd1 vssd1 vccd1 vccd1 _8487_/A sky130_fd_sc_hd__xnor2_1
X_5663_ _5974_/A _5659_/Y _6063_/A vssd1 vssd1 vccd1 vccd1 _5706_/A sky130_fd_sc_hd__a21oi_2
XFILLER_30_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8382_ _8382_/A _8385_/B vssd1 vssd1 vccd1 vccd1 _8445_/C sky130_fd_sc_hd__nand2_1
X_7402_ _7402_/A _7402_/B vssd1 vssd1 vccd1 vccd1 _7422_/A sky130_fd_sc_hd__xnor2_1
X_4614_ _8580_/Q _4614_/B vssd1 vssd1 vccd1 vccd1 _4619_/C sky130_fd_sc_hd__and2_1
X_5594_ _5795_/A vssd1 vssd1 vccd1 vccd1 _5742_/A sky130_fd_sc_hd__buf_2
X_7333_ _7333_/A _7333_/B _7333_/C vssd1 vssd1 vccd1 vccd1 _7333_/Y sky130_fd_sc_hd__nor3_2
X_4545_ _4545_/A vssd1 vssd1 vccd1 vccd1 _8866_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_89_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7264_ _7264_/A _7264_/B vssd1 vssd1 vccd1 vccd1 _7313_/B sky130_fd_sc_hd__xnor2_2
XFILLER_89_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4476_ _5226_/B _4705_/A _4662_/A vssd1 vssd1 vccd1 vccd1 _4709_/A sky130_fd_sc_hd__and3_1
X_7195_ _7195_/A _7195_/B vssd1 vssd1 vccd1 vccd1 _7289_/B sky130_fd_sc_hd__xnor2_2
X_6215_ _6215_/A _6215_/B _6215_/C vssd1 vssd1 vccd1 vccd1 _6217_/A sky130_fd_sc_hd__or3_1
XFILLER_85_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6146_ _6322_/A _6322_/B _6327_/B vssd1 vssd1 vccd1 vccd1 _6302_/B sky130_fd_sc_hd__and3_1
XFILLER_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6077_ _6077_/A _6077_/B vssd1 vssd1 vccd1 vccd1 _6087_/A sky130_fd_sc_hd__xnor2_1
X_5028_ _5176_/A _5151_/A _5118_/D vssd1 vssd1 vccd1 vccd1 _5028_/X sky130_fd_sc_hd__or3_1
XFILLER_26_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6979_ _6979_/A _6979_/B vssd1 vssd1 vccd1 vccd1 _6980_/B sky130_fd_sc_hd__xnor2_1
XFILLER_41_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8718_ input3/X _8718_/D vssd1 vssd1 vccd1 vccd1 _8718_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8649_ input3/X _8649_/D vssd1 vssd1 vccd1 vccd1 _8649_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8803__81 vssd1 vssd1 vccd1 vccd1 _8803__81/HI _8912_/A sky130_fd_sc_hd__conb_1
XFILLER_63_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4330_ _4333_/A vssd1 vssd1 vccd1 vccd1 _4330_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6000_ _6000_/A _6000_/B vssd1 vssd1 vccd1 vccd1 _6207_/B sky130_fd_sc_hd__nand2_1
XFILLER_79_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7951_ _7894_/B _7894_/C _7894_/A vssd1 vssd1 vccd1 vccd1 _7978_/A sky130_fd_sc_hd__a21bo_1
XFILLER_82_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7882_ _7882_/A _7882_/B _7882_/C vssd1 vssd1 vccd1 vccd1 _7894_/A sky130_fd_sc_hd__nand3_1
X_6902_ _6919_/A _6919_/B vssd1 vssd1 vccd1 vccd1 _7045_/B sky130_fd_sc_hd__or2_1
XFILLER_54_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6833_ _6833_/A _6833_/B vssd1 vssd1 vccd1 vccd1 _6834_/B sky130_fd_sc_hd__xnor2_1
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6764_ _6719_/A _6763_/Y _6689_/X vssd1 vssd1 vccd1 vccd1 _6766_/A sky130_fd_sc_hd__a21oi_2
XFILLER_50_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8503_ _8503_/A _8503_/B _8503_/C vssd1 vssd1 vccd1 vccd1 _8503_/X sky130_fd_sc_hd__and3_1
X_6695_ _6695_/A vssd1 vssd1 vccd1 vccd1 _7293_/B sky130_fd_sc_hd__clkbuf_2
X_5715_ _5602_/A _5715_/B vssd1 vssd1 vccd1 vccd1 _5715_/X sky130_fd_sc_hd__and2b_1
X_8434_ _8427_/A _8432_/B _8427_/B vssd1 vssd1 vccd1 vccd1 _8490_/B sky130_fd_sc_hd__a21bo_1
X_5646_ _5646_/A _5832_/A vssd1 vssd1 vccd1 vccd1 _6053_/A sky130_fd_sc_hd__nand2_1
X_8365_ _8365_/A _8365_/B vssd1 vssd1 vccd1 vccd1 _8366_/B sky130_fd_sc_hd__xor2_1
X_5577_ _5554_/A _5577_/B vssd1 vssd1 vccd1 vccd1 _5718_/A sky130_fd_sc_hd__nand2b_1
X_8296_ _8296_/A _8296_/B vssd1 vssd1 vccd1 vccd1 _8353_/B sky130_fd_sc_hd__xnor2_1
X_7316_ _7301_/A _7301_/B _7315_/X vssd1 vssd1 vccd1 vccd1 _7323_/A sky130_fd_sc_hd__a21o_1
X_4528_ _5180_/A vssd1 vssd1 vccd1 vccd1 _5083_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7247_ _7296_/C _7248_/B _7246_/X vssd1 vssd1 vccd1 vccd1 _7264_/A sky130_fd_sc_hd__a21o_2
XFILLER_49_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4459_ _4459_/A vssd1 vssd1 vccd1 vccd1 _4459_/Y sky130_fd_sc_hd__inv_2
X_7178_ _6697_/A _7299_/A _7315_/A _7251_/B vssd1 vssd1 vccd1 vccd1 _7239_/B sky130_fd_sc_hd__a22o_1
XFILLER_58_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6129_ _5800_/A _6083_/C _6145_/A vssd1 vssd1 vccd1 vccd1 _6131_/B sky130_fd_sc_hd__o21ba_1
XFILLER_100_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5500_ _8600_/Q vssd1 vssd1 vccd1 vccd1 _6608_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6480_ _7525_/A vssd1 vssd1 vccd1 vccd1 _7537_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5431_ _5428_/A _5419_/X _5429_/X _5430_/Y _4743_/X vssd1 vssd1 vccd1 vccd1 _8650_/D
+ sky130_fd_sc_hd__o221a_1
X_8150_ _8146_/B _8149_/B _8149_/Y vssd1 vssd1 vccd1 vccd1 _8151_/B sky130_fd_sc_hd__o21ai_1
X_5362_ _5366_/C _5362_/B vssd1 vssd1 vccd1 vccd1 _8638_/D sky130_fd_sc_hd__nor2_1
X_8081_ _8256_/A _8081_/B vssd1 vssd1 vccd1 vccd1 _8083_/B sky130_fd_sc_hd__nor2_1
X_7101_ _7115_/B _7101_/B _7101_/C _7101_/D vssd1 vssd1 vccd1 vccd1 _7103_/A sky130_fd_sc_hd__nand4_1
XFILLER_99_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7032_ _7032_/A _7032_/B vssd1 vssd1 vccd1 vccd1 _7034_/B sky130_fd_sc_hd__xor2_1
X_5293_ _8620_/Q _5300_/B vssd1 vssd1 vccd1 vccd1 _5293_/X sky130_fd_sc_hd__or2_1
XFILLER_67_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7934_ _7817_/X _8056_/B _7800_/B _7933_/X vssd1 vssd1 vccd1 vccd1 _7936_/B sky130_fd_sc_hd__a31oi_1
XFILLER_35_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7865_ _7889_/A _7865_/B _7865_/C vssd1 vssd1 vccd1 vccd1 _7867_/B sky130_fd_sc_hd__or3_1
XFILLER_70_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8794__72 vssd1 vssd1 vccd1 vccd1 _8794__72/HI _8903_/A sky130_fd_sc_hd__conb_1
XFILLER_51_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6816_ _6685_/A _6763_/Y _6689_/X _6815_/X vssd1 vssd1 vccd1 vccd1 _6949_/A sky130_fd_sc_hd__a211o_2
X_7796_ _7796_/A _7796_/B vssd1 vssd1 vccd1 vccd1 _7796_/X sky130_fd_sc_hd__or2_1
X_6747_ _7226_/B _7236_/B _7265_/B vssd1 vssd1 vccd1 vccd1 _6748_/B sky130_fd_sc_hd__o21ai_1
XFILLER_11_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6678_ _7177_/A vssd1 vssd1 vccd1 vccd1 _7297_/B sky130_fd_sc_hd__clkbuf_2
X_8417_ _8417_/A _8417_/B vssd1 vssd1 vccd1 vccd1 _8418_/B sky130_fd_sc_hd__xor2_2
X_5629_ _5660_/A _5629_/B vssd1 vssd1 vccd1 vccd1 _5646_/A sky130_fd_sc_hd__xnor2_1
X_8348_ _8351_/B _8348_/B vssd1 vssd1 vccd1 vccd1 _8352_/B sky130_fd_sc_hd__xnor2_1
XFILLER_2_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8279_ _8301_/B _8279_/B vssd1 vssd1 vccd1 vccd1 _8288_/A sky130_fd_sc_hd__nand2_1
XFILLER_2_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5980_ _5980_/A _6284_/S vssd1 vssd1 vccd1 vccd1 _5980_/X sky130_fd_sc_hd__or2_1
X_4931_ _5098_/D _4976_/C vssd1 vssd1 vccd1 vccd1 _5175_/B sky130_fd_sc_hd__nor2_2
XFILLER_17_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7650_ _7912_/A vssd1 vssd1 vccd1 vccd1 _7790_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_60_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4862_ _5087_/A _5119_/C vssd1 vssd1 vccd1 vccd1 _5072_/B sky130_fd_sc_hd__or2_2
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6601_ _6608_/B _8704_/Q vssd1 vssd1 vccd1 vccd1 _6836_/A sky130_fd_sc_hd__or2b_1
XFILLER_60_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7581_ _8564_/A vssd1 vssd1 vccd1 vccd1 _7581_/X sky130_fd_sc_hd__buf_2
X_4793_ _4535_/C _4795_/B _4820_/A vssd1 vssd1 vccd1 vccd1 _4794_/B sky130_fd_sc_hd__o21bai_1
X_6532_ _6527_/B _6529_/B _6525_/Y vssd1 vssd1 vccd1 vccd1 _6533_/C sky130_fd_sc_hd__a21oi_1
X_6463_ _8683_/Q _6463_/B vssd1 vssd1 vccd1 vccd1 _6465_/A sky130_fd_sc_hd__and2_1
X_8202_ _8202_/A _8202_/B vssd1 vssd1 vccd1 vccd1 _8241_/A sky130_fd_sc_hd__xor2_1
X_5414_ _5414_/A _8646_/Q vssd1 vssd1 vccd1 vccd1 _5416_/B sky130_fd_sc_hd__xor2_1
X_8133_ _8133_/A _8203_/B vssd1 vssd1 vccd1 vccd1 _8138_/A sky130_fd_sc_hd__xnor2_2
X_6394_ _8666_/Q _8665_/Q vssd1 vssd1 vccd1 vccd1 _6400_/A sky130_fd_sc_hd__nor2_1
XFILLER_99_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5345_ _5345_/A vssd1 vssd1 vccd1 vccd1 _8633_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8064_ _8371_/A _8363_/A vssd1 vssd1 vccd1 vccd1 _8437_/A sky130_fd_sc_hd__xnor2_2
X_5276_ _8655_/Q _5271_/X _5275_/X _5273_/X vssd1 vssd1 vccd1 vccd1 _8613_/D sky130_fd_sc_hd__o211a_1
X_7015_ _7149_/B _7015_/B vssd1 vssd1 vccd1 vccd1 _7016_/B sky130_fd_sc_hd__xnor2_2
XFILLER_68_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7917_ _7998_/A _7998_/B vssd1 vssd1 vccd1 vccd1 _7923_/A sky130_fd_sc_hd__xnor2_1
X_8897_ _8897_/A _4408_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[6] sky130_fd_sc_hd__ebufn_8
X_7848_ _7848_/A _8512_/A vssd1 vssd1 vccd1 vccd1 _7849_/B sky130_fd_sc_hd__or2_1
XFILLER_11_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7779_ _7779_/A vssd1 vssd1 vccd1 vccd1 _8283_/A sky130_fd_sc_hd__inv_2
XFILLER_51_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5130_ _5130_/A _5130_/B vssd1 vssd1 vccd1 vccd1 _5137_/C sky130_fd_sc_hd__or2_1
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5061_ _5091_/A vssd1 vssd1 vccd1 vccd1 _5214_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_65_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5963_ _5964_/B _6182_/A _5922_/A vssd1 vssd1 vccd1 vccd1 _5965_/B sky130_fd_sc_hd__a21o_1
XFILLER_18_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8764__42 vssd1 vssd1 vccd1 vccd1 _8764__42/HI _8859_/A sky130_fd_sc_hd__conb_1
X_7702_ _8722_/Q vssd1 vssd1 vccd1 vccd1 _7702_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4914_ _4887_/X _4907_/X _4728_/A _5238_/A vssd1 vssd1 vccd1 vccd1 _4914_/X sky130_fd_sc_hd__a211o_1
XFILLER_80_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8682_ input3/X _8682_/D vssd1 vssd1 vccd1 vccd1 _8682_/Q sky130_fd_sc_hd__dfxtp_1
X_5894_ _6007_/A _5726_/A _5809_/A _5809_/B vssd1 vssd1 vccd1 vccd1 _5902_/A sky130_fd_sc_hd__a22o_1
X_4845_ _4859_/A vssd1 vssd1 vccd1 vccd1 _5041_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7633_ _8710_/Q _8607_/Q vssd1 vssd1 vccd1 vccd1 _7633_/X sky130_fd_sc_hd__and2b_1
X_7564_ _7616_/B vssd1 vssd1 vccd1 vccd1 _7615_/B sky130_fd_sc_hd__clkbuf_2
X_4776_ _7547_/A _4776_/B _4778_/B vssd1 vssd1 vccd1 vccd1 _4777_/A sky130_fd_sc_hd__and3_1
X_6515_ _6567_/A _6516_/B vssd1 vssd1 vccd1 vccd1 _6515_/Y sky130_fd_sc_hd__nor2_1
X_7495_ _7495_/A _7495_/B vssd1 vssd1 vccd1 vccd1 _7496_/B sky130_fd_sc_hd__and2_1
X_6446_ _8677_/Q _6445_/B _6419_/X vssd1 vssd1 vccd1 vccd1 _6447_/B sky130_fd_sc_hd__o21ai_1
X_6377_ _5419_/X _6376_/X _8664_/Q vssd1 vssd1 vccd1 vccd1 _6379_/A sky130_fd_sc_hd__a21oi_1
XFILLER_102_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8116_ _8326_/B _8116_/B _8116_/C vssd1 vssd1 vccd1 vccd1 _8230_/A sky130_fd_sc_hd__and3b_1
X_5328_ _6475_/B _5330_/C _5374_/A vssd1 vssd1 vccd1 vccd1 _5328_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8047_ _8047_/A _8047_/B vssd1 vssd1 vccd1 vccd1 _8103_/B sky130_fd_sc_hd__xor2_2
XFILLER_75_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5259_ _5259_/A _5259_/B _5259_/C vssd1 vssd1 vccd1 vccd1 _5259_/X sky130_fd_sc_hd__or3_1
XFILLER_28_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4630_ _4632_/B _4639_/B _4630_/C vssd1 vssd1 vccd1 vccd1 _4631_/A sky130_fd_sc_hd__and3b_1
XFILLER_8_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4561_ _8616_/Q _4563_/B vssd1 vssd1 vccd1 vccd1 _4562_/A sky130_fd_sc_hd__and2_1
XFILLER_8_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6300_ _6300_/A _6300_/B vssd1 vssd1 vccd1 vccd1 _6301_/B sky130_fd_sc_hd__nand2_1
X_7280_ _7279_/B _7280_/B vssd1 vssd1 vccd1 vccd1 _7280_/X sky130_fd_sc_hd__and2b_1
X_4492_ _7634_/A vssd1 vssd1 vccd1 vccd1 _5620_/A sky130_fd_sc_hd__buf_2
X_6231_ _6231_/A _6231_/B vssd1 vssd1 vccd1 vccd1 _6232_/B sky130_fd_sc_hd__nor2_1
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6162_ _6311_/A _6311_/B vssd1 vssd1 vccd1 vccd1 _6312_/A sky130_fd_sc_hd__nand2_1
XFILLER_97_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5113_ _5113_/A _5113_/B vssd1 vssd1 vccd1 vccd1 _5113_/Y sky130_fd_sc_hd__nand2_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6093_ _6060_/B _6091_/X _6090_/Y _6084_/X vssd1 vssd1 vccd1 vccd1 _6095_/B sky130_fd_sc_hd__o211a_1
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5044_ _5253_/C _5172_/C _5118_/D _5044_/D vssd1 vssd1 vccd1 vccd1 _5044_/X sky130_fd_sc_hd__or4_1
XFILLER_38_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6995_ _6995_/A _6995_/B vssd1 vssd1 vccd1 vccd1 _7087_/A sky130_fd_sc_hd__nor2_1
XFILLER_80_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5946_ _5946_/A _5946_/B vssd1 vssd1 vccd1 vccd1 _5946_/Y sky130_fd_sc_hd__nor2_1
X_5877_ _5815_/A _5877_/B vssd1 vssd1 vccd1 vccd1 _5877_/X sky130_fd_sc_hd__and2b_1
XFILLER_21_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8665_ input3/X _8665_/D vssd1 vssd1 vccd1 vccd1 _8665_/Q sky130_fd_sc_hd__dfxtp_1
X_7616_ _7616_/A _7616_/B vssd1 vssd1 vccd1 vccd1 _7621_/B sky130_fd_sc_hd__or2_1
X_4828_ _4872_/C _4828_/B vssd1 vssd1 vccd1 vccd1 _5109_/B sky130_fd_sc_hd__nor2_2
X_8596_ input3/X _8596_/D vssd1 vssd1 vccd1 vccd1 _8596_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_5_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4759_ _5290_/A _4856_/A _4495_/A vssd1 vssd1 vccd1 vccd1 _4761_/B sky130_fd_sc_hd__o21bai_1
X_7547_ _7547_/A _7547_/B _7547_/C vssd1 vssd1 vccd1 vccd1 _7548_/A sky130_fd_sc_hd__and3_1
X_7478_ _7478_/A _7480_/B vssd1 vssd1 vccd1 vccd1 _7479_/B sky130_fd_sc_hd__nand2_1
X_6429_ _6429_/A _6429_/B vssd1 vssd1 vccd1 vccd1 _8671_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6780_ _7194_/B vssd1 vssd1 vccd1 vccd1 _6869_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_62_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5800_ _5800_/A _6213_/B vssd1 vssd1 vccd1 vccd1 _5800_/X sky130_fd_sc_hd__or2_1
X_8734__12 vssd1 vssd1 vccd1 vccd1 _8734__12/HI _8829_/A sky130_fd_sc_hd__conb_1
XFILLER_62_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5731_ _5731_/A vssd1 vssd1 vccd1 vccd1 _5803_/B sky130_fd_sc_hd__buf_2
X_8450_ _8441_/X _8442_/Y _8448_/Y _8449_/Y vssd1 vssd1 vccd1 vccd1 _8451_/B sky130_fd_sc_hd__a31o_1
X_5662_ _5660_/Y _5629_/B _5658_/A _5923_/B vssd1 vssd1 vccd1 vccd1 _6063_/A sky130_fd_sc_hd__o211a_2
X_8381_ _8381_/A _8323_/B vssd1 vssd1 vccd1 vccd1 _8388_/B sky130_fd_sc_hd__or2b_1
X_7401_ _7296_/A _7296_/C _7400_/X vssd1 vssd1 vccd1 vccd1 _7402_/B sky130_fd_sc_hd__a21oi_2
X_4613_ _4613_/A vssd1 vssd1 vccd1 vccd1 _8579_/D sky130_fd_sc_hd__clkbuf_1
X_5593_ _5551_/A _5895_/A _5553_/B _5553_/A vssd1 vssd1 vccd1 vccd1 _5740_/A sky130_fd_sc_hd__a22o_1
X_7332_ _7332_/A _7332_/B vssd1 vssd1 vccd1 vccd1 _7333_/C sky130_fd_sc_hd__xnor2_1
X_4544_ _8612_/Q _4552_/B vssd1 vssd1 vccd1 vccd1 _4545_/A sky130_fd_sc_hd__and2_1
X_7263_ _7262_/B _7262_/C _7262_/A vssd1 vssd1 vccd1 vccd1 _7334_/C sky130_fd_sc_hd__a21o_1
X_6214_ _6214_/A _6214_/B vssd1 vssd1 vccd1 vccd1 _6215_/C sky130_fd_sc_hd__nor2_1
X_4475_ _7753_/A _7688_/B _4475_/C _4723_/A vssd1 vssd1 vccd1 vccd1 _4520_/A sky130_fd_sc_hd__or4b_1
X_7194_ _7223_/A _7194_/B vssd1 vssd1 vccd1 vccd1 _7195_/B sky130_fd_sc_hd__nor2_1
X_6145_ _6145_/A _6145_/B vssd1 vssd1 vccd1 vccd1 _6327_/B sky130_fd_sc_hd__nor2_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6076_ _6167_/A _6307_/B vssd1 vssd1 vccd1 vccd1 _6076_/Y sky130_fd_sc_hd__xnor2_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5027_ _5185_/C _5027_/B vssd1 vssd1 vccd1 vccd1 _5118_/D sky130_fd_sc_hd__or2_2
XFILLER_80_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6978_ _6978_/A _6978_/B vssd1 vssd1 vccd1 vccd1 _6979_/B sky130_fd_sc_hd__xnor2_2
X_8717_ input3/X _8717_/D vssd1 vssd1 vccd1 vccd1 _8717_/Q sky130_fd_sc_hd__dfxtp_1
X_5929_ _5950_/A _5929_/B vssd1 vssd1 vccd1 vccd1 _5932_/A sky130_fd_sc_hd__xor2_1
XFILLER_41_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8648_ input3/X _8648_/D vssd1 vssd1 vccd1 vccd1 _8648_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8579_ input3/X _8579_/D vssd1 vssd1 vccd1 vccd1 _8579_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7950_ _8207_/A _8331_/A _7898_/D _7949_/X vssd1 vssd1 vccd1 vccd1 _7982_/A sky130_fd_sc_hd__a31o_1
XFILLER_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7881_ _7880_/A _7880_/B _7880_/C vssd1 vssd1 vccd1 vccd1 _7882_/C sky130_fd_sc_hd__a21o_1
X_6901_ _7296_/B _7246_/B vssd1 vssd1 vccd1 vccd1 _7045_/A sky130_fd_sc_hd__nand2_1
X_6832_ _6951_/A _7023_/A vssd1 vssd1 vccd1 vccd1 _6833_/B sky130_fd_sc_hd__xor2_1
X_6763_ _7237_/B _7177_/A _7237_/C _6718_/S vssd1 vssd1 vccd1 vccd1 _6763_/Y sky130_fd_sc_hd__o31ai_2
X_8502_ _8502_/A _8502_/B vssd1 vssd1 vccd1 vccd1 _8502_/Y sky130_fd_sc_hd__xnor2_1
X_6694_ _6798_/B _7048_/C vssd1 vssd1 vccd1 vccd1 _6723_/A sky130_fd_sc_hd__nor2_1
X_5714_ _6061_/A _6061_/B _5713_/Y vssd1 vssd1 vccd1 vccd1 _5771_/A sky130_fd_sc_hd__a21boi_1
X_8433_ _8492_/B _8492_/C _8493_/B _8492_/A vssd1 vssd1 vccd1 vccd1 _8490_/A sky130_fd_sc_hd__a211o_1
X_5645_ _5657_/A _5645_/B vssd1 vssd1 vccd1 vccd1 _5832_/A sky130_fd_sc_hd__nand2_1
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8364_ _8364_/A _8443_/B vssd1 vssd1 vccd1 vccd1 _8365_/B sky130_fd_sc_hd__xnor2_1
X_5576_ _5569_/A _5576_/B vssd1 vssd1 vccd1 vccd1 _5602_/A sky130_fd_sc_hd__and2b_1
XFILLER_104_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8295_ _8295_/A _8295_/B vssd1 vssd1 vccd1 vccd1 _8296_/B sky130_fd_sc_hd__xnor2_1
X_7315_ _7315_/A _7418_/C _7315_/C vssd1 vssd1 vccd1 vccd1 _7315_/X sky130_fd_sc_hd__and3_1
XFILLER_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4527_ _8592_/Q vssd1 vssd1 vccd1 vccd1 _5180_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4458_ _4459_/A vssd1 vssd1 vccd1 vccd1 _4458_/Y sky130_fd_sc_hd__inv_2
X_7246_ _7293_/A _7246_/B _7294_/A vssd1 vssd1 vccd1 vccd1 _7246_/X sky130_fd_sc_hd__and3_1
XFILLER_49_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7177_ _7177_/A _7243_/A vssd1 vssd1 vccd1 vccd1 _7251_/B sky130_fd_sc_hd__xnor2_2
X_4389_ _4389_/A vssd1 vssd1 vccd1 vccd1 _4389_/Y sky130_fd_sc_hd__inv_2
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6128_ _6142_/A _6128_/B _6128_/C vssd1 vssd1 vccd1 vccd1 _6145_/A sky130_fd_sc_hd__and3_1
XFILLER_100_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6059_ _6060_/A _6059_/B _6058_/X vssd1 vssd1 vccd1 vccd1 _6060_/B sky130_fd_sc_hd__nor3b_1
XFILLER_45_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5430_ _5422_/A _5424_/Y _5428_/X _5419_/A vssd1 vssd1 vccd1 vccd1 _5430_/Y sky130_fd_sc_hd__o31ai_1
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5361_ _8638_/Q _5359_/A _5357_/X vssd1 vssd1 vccd1 vccd1 _5362_/B sky130_fd_sc_hd__o21ai_1
X_8080_ _8079_/A _8079_/B _8079_/C vssd1 vssd1 vccd1 vccd1 _8081_/B sky130_fd_sc_hd__a21oi_1
X_7100_ _7100_/A _7100_/B vssd1 vssd1 vccd1 vccd1 _7106_/A sky130_fd_sc_hd__xnor2_1
X_5292_ _8718_/Q _5285_/X _5291_/X _5283_/X vssd1 vssd1 vccd1 vccd1 _8619_/D sky130_fd_sc_hd__o211a_1
X_7031_ _6744_/A _7265_/B _7031_/S vssd1 vssd1 vccd1 vccd1 _7032_/B sky130_fd_sc_hd__mux2_1
XFILLER_28_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7933_ _7902_/A _7933_/B vssd1 vssd1 vccd1 vccd1 _7933_/X sky130_fd_sc_hd__and2b_1
XFILLER_55_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7864_ _7864_/A _7864_/B _7877_/A vssd1 vssd1 vccd1 vccd1 _7865_/C sky130_fd_sc_hd__and3_1
XFILLER_63_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6815_ _6717_/X _6815_/B _6815_/C vssd1 vssd1 vccd1 vccd1 _6815_/X sky130_fd_sc_hd__and3b_1
X_7795_ _7924_/A _7924_/B vssd1 vssd1 vccd1 vccd1 _7801_/A sky130_fd_sc_hd__xor2_1
X_6746_ _6842_/A vssd1 vssd1 vccd1 vccd1 _7265_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6677_ _7249_/B _6700_/B _6769_/A vssd1 vssd1 vccd1 vccd1 _6724_/A sky130_fd_sc_hd__nand3_1
X_8416_ _8416_/A _8416_/B vssd1 vssd1 vccd1 vccd1 _8417_/B sky130_fd_sc_hd__nor2_1
X_5628_ _5617_/X _5642_/A _5631_/B _5633_/B vssd1 vssd1 vccd1 vccd1 _5629_/B sky130_fd_sc_hd__a31o_1
X_8347_ _8347_/A _8347_/B vssd1 vssd1 vccd1 vccd1 _8348_/B sky130_fd_sc_hd__xnor2_1
X_5559_ _5879_/A _5559_/B _5595_/A vssd1 vssd1 vccd1 vccd1 _5567_/A sky130_fd_sc_hd__and3_1
XFILLER_78_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8278_ _7666_/A _7671_/A _8508_/A vssd1 vssd1 vccd1 vccd1 _8279_/B sky130_fd_sc_hd__a21o_1
XFILLER_104_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7229_ _7229_/A _7229_/B vssd1 vssd1 vccd1 vccd1 _7376_/A sky130_fd_sc_hd__xnor2_1
XFILLER_76_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4930_ _4930_/A _4930_/B vssd1 vssd1 vccd1 vccd1 _4976_/C sky130_fd_sc_hd__nor2_1
XFILLER_24_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4861_ _4861_/A _4865_/B vssd1 vssd1 vccd1 vccd1 _5119_/C sky130_fd_sc_hd__nor2_1
X_6600_ _6635_/A _6600_/B vssd1 vssd1 vccd1 vccd1 _6737_/A sky130_fd_sc_hd__nor2_2
X_7580_ _8535_/S vssd1 vssd1 vccd1 vccd1 _8564_/A sky130_fd_sc_hd__clkbuf_2
X_4792_ _5620_/A _4795_/B _4820_/A vssd1 vssd1 vccd1 vccd1 _4848_/B sky130_fd_sc_hd__or3b_1
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6531_ _6536_/A _6531_/B vssd1 vssd1 vccd1 vccd1 _6540_/A sky130_fd_sc_hd__nand2_1
XFILLER_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6462_ _6462_/A vssd1 vssd1 vccd1 vccd1 _8682_/D sky130_fd_sc_hd__clkbuf_1
X_8201_ _8201_/A _8201_/B vssd1 vssd1 vccd1 vccd1 _8202_/B sky130_fd_sc_hd__xnor2_1
X_5413_ _5413_/A vssd1 vssd1 vccd1 vccd1 _5413_/X sky130_fd_sc_hd__buf_2
X_6393_ _8685_/Q _6393_/B vssd1 vssd1 vccd1 vccd1 _6406_/B sky130_fd_sc_hd__nand2_1
XFILLER_99_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8132_ _8132_/A _8132_/B vssd1 vssd1 vccd1 vccd1 _8203_/B sky130_fd_sc_hd__xnor2_2
X_5344_ _5346_/B _5344_/B _5354_/B vssd1 vssd1 vccd1 vccd1 _5345_/A sky130_fd_sc_hd__and3b_1
XFILLER_99_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8063_ _8063_/A vssd1 vssd1 vccd1 vccd1 _8371_/A sky130_fd_sc_hd__buf_2
X_5275_ _8613_/Q _5275_/B vssd1 vssd1 vccd1 vccd1 _5275_/X sky130_fd_sc_hd__or2_1
X_7014_ _6982_/A _6982_/B _7013_/Y vssd1 vssd1 vccd1 vccd1 _7015_/B sky130_fd_sc_hd__o21a_1
XFILLER_87_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7916_ _7916_/A _7984_/B vssd1 vssd1 vccd1 vccd1 _7998_/B sky130_fd_sc_hd__xnor2_1
X_8896_ _8896_/A _4410_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[5] sky130_fd_sc_hd__ebufn_8
XFILLER_36_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7847_ _7847_/A vssd1 vssd1 vccd1 vccd1 _7847_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7778_ _7850_/A _7850_/B vssd1 vssd1 vccd1 vccd1 _7807_/A sky130_fd_sc_hd__xnor2_1
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6729_ _6900_/A _6729_/B vssd1 vssd1 vccd1 vccd1 _6730_/B sky130_fd_sc_hd__xnor2_1
XFILLER_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5060_ _5060_/A _5190_/C _5060_/C _5059_/X vssd1 vssd1 vccd1 vccd1 _5060_/X sky130_fd_sc_hd__or4b_1
XFILLER_84_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5962_ _5962_/A _6107_/B vssd1 vssd1 vccd1 vccd1 _6182_/A sky130_fd_sc_hd__or2_1
XFILLER_18_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7701_ _7701_/A _7701_/B vssd1 vssd1 vccd1 vccd1 _7717_/B sky130_fd_sc_hd__nor2_1
XFILLER_52_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4913_ _5241_/A vssd1 vssd1 vccd1 vccd1 _5238_/A sky130_fd_sc_hd__clkbuf_2
X_5893_ _5897_/B vssd1 vssd1 vccd1 vccd1 _6007_/A sky130_fd_sc_hd__clkbuf_2
X_8681_ input3/X _8681_/D vssd1 vssd1 vccd1 vccd1 _8681_/Q sky130_fd_sc_hd__dfxtp_1
X_7632_ _7649_/A _7654_/B _7631_/X vssd1 vssd1 vccd1 vccd1 _7636_/A sky130_fd_sc_hd__a21oi_1
X_4844_ _5015_/A _4933_/A _5245_/C vssd1 vssd1 vccd1 vccd1 _5042_/A sky130_fd_sc_hd__or3_1
XFILLER_33_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7563_ _8707_/Q vssd1 vssd1 vccd1 vccd1 _7616_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4775_ _4775_/A _5263_/A _4775_/C vssd1 vssd1 vccd1 vccd1 _4778_/B sky130_fd_sc_hd__nand3_1
XFILLER_20_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6514_ _6514_/A _8687_/Q vssd1 vssd1 vccd1 vccd1 _6516_/B sky130_fd_sc_hd__xor2_1
X_7494_ _7494_/A vssd1 vssd1 vccd1 vccd1 _7494_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6445_ _8677_/Q _6445_/B vssd1 vssd1 vccd1 vccd1 _6450_/C sky130_fd_sc_hd__and2_1
X_6376_ _6372_/A _6375_/X _6376_/S vssd1 vssd1 vccd1 vccd1 _6376_/X sky130_fd_sc_hd__mux2_1
X_8115_ _8115_/A vssd1 vssd1 vccd1 vccd1 _8326_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_5327_ _5330_/C _5327_/B vssd1 vssd1 vccd1 vccd1 _8627_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8046_ _8031_/A _8043_/Y _8158_/A vssd1 vssd1 vccd1 vccd1 _8047_/B sky130_fd_sc_hd__a21oi_2
XFILLER_87_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5258_ _5243_/C _5252_/X _5253_/X _5257_/X _5248_/B vssd1 vssd1 vccd1 vccd1 _5259_/C
+ sky130_fd_sc_hd__o32a_1
XFILLER_68_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5189_ _5040_/A _5029_/B _5184_/X _5185_/X _5188_/X vssd1 vssd1 vccd1 vccd1 _5190_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_83_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8879_ _8879_/A _4398_/Y vssd1 vssd1 vccd1 vccd1 io_out[26] sky130_fd_sc_hd__ebufn_8
XFILLER_12_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4560_ _4560_/A vssd1 vssd1 vccd1 vccd1 _8877_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_8_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4491_ _8607_/Q vssd1 vssd1 vccd1 vccd1 _7634_/A sky130_fd_sc_hd__clkbuf_4
X_6230_ _6231_/A _6230_/B _6230_/C vssd1 vssd1 vccd1 vccd1 _6232_/A sky130_fd_sc_hd__and3_1
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6161_ _6161_/A _6161_/B vssd1 vssd1 vccd1 vccd1 _6311_/B sky130_fd_sc_hd__xor2_1
XFILLER_97_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5112_ _5106_/X _5107_/X _5111_/X vssd1 vssd1 vccd1 vccd1 _5113_/B sky130_fd_sc_hd__o21ai_1
XFILLER_97_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6092_ _6084_/X _6090_/Y _6091_/X _6060_/B vssd1 vssd1 vccd1 vccd1 _6096_/A sky130_fd_sc_hd__a211oi_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5043_ _5180_/A _5245_/D _5046_/B vssd1 vssd1 vccd1 vccd1 _5044_/D sky130_fd_sc_hd__or3_1
XFILLER_65_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6994_ _6991_/X _6992_/X _6995_/A _6993_/Y vssd1 vssd1 vccd1 vccd1 _6995_/B sky130_fd_sc_hd__a211oi_2
XFILLER_92_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5945_ _5937_/A _5937_/B _5938_/A _5936_/A vssd1 vssd1 vccd1 vccd1 _6027_/A sky130_fd_sc_hd__a31o_1
X_5876_ _5920_/B _5876_/B vssd1 vssd1 vccd1 vccd1 _5918_/A sky130_fd_sc_hd__xor2_1
XFILLER_33_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8664_ input3/X _8664_/D vssd1 vssd1 vccd1 vccd1 _8664_/Q sky130_fd_sc_hd__dfxtp_1
X_7615_ _7616_/A _7615_/B vssd1 vssd1 vccd1 vccd1 _7617_/A sky130_fd_sc_hd__nand2_1
X_4827_ _4822_/C _4872_/B _4848_/A vssd1 vssd1 vccd1 vccd1 _4828_/B sky130_fd_sc_hd__a21oi_1
X_8595_ input3/X _8595_/D vssd1 vssd1 vccd1 vccd1 _8595_/Q sky130_fd_sc_hd__dfxtp_2
X_7546_ _7540_/A _7545_/C _7545_/A vssd1 vssd1 vccd1 vccd1 _7547_/C sky130_fd_sc_hd__o21ai_1
X_4758_ _4758_/A vssd1 vssd1 vccd1 vccd1 _8605_/D sky130_fd_sc_hd__clkbuf_1
X_7477_ _7477_/A _7477_/B vssd1 vssd1 vccd1 vccd1 _7479_/A sky130_fd_sc_hd__nand2_1
X_4689_ _4695_/A _4688_/X _4717_/A vssd1 vssd1 vccd1 vccd1 _8594_/D sky130_fd_sc_hd__a21boi_1
X_6428_ _6430_/A _6430_/C _6427_/X vssd1 vssd1 vccd1 vccd1 _6429_/B sky130_fd_sc_hd__o21ai_1
X_6359_ _6352_/B _6354_/B _6352_/A vssd1 vssd1 vccd1 vccd1 _6359_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_102_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8029_ _8117_/S _8029_/B vssd1 vssd1 vccd1 vccd1 _8109_/A sky130_fd_sc_hd__xnor2_2
XFILLER_88_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5730_ _5789_/A _5789_/B vssd1 vssd1 vccd1 vccd1 _5738_/A sky130_fd_sc_hd__xnor2_2
XFILLER_50_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7400_ _7297_/A _7378_/B _7418_/C _6647_/A vssd1 vssd1 vccd1 vccd1 _7400_/X sky130_fd_sc_hd__o22a_1
X_5661_ _6042_/A _5957_/B vssd1 vssd1 vccd1 vccd1 _5923_/B sky130_fd_sc_hd__nor2_2
X_8380_ _8380_/A _8322_/A vssd1 vssd1 vccd1 vccd1 _8388_/A sky130_fd_sc_hd__or2b_1
X_4612_ _4614_/B _4639_/B _4612_/C vssd1 vssd1 vccd1 vccd1 _4613_/A sky130_fd_sc_hd__and3b_1
X_5592_ _6003_/A vssd1 vssd1 vccd1 vccd1 _5895_/A sky130_fd_sc_hd__clkbuf_2
X_7331_ _7330_/A _7330_/C _7330_/B vssd1 vssd1 vccd1 vccd1 _7333_/B sky130_fd_sc_hd__a21oi_1
X_4543_ _4567_/B vssd1 vssd1 vccd1 vccd1 _4552_/B sky130_fd_sc_hd__clkbuf_2
X_7262_ _7262_/A _7262_/B _7262_/C vssd1 vssd1 vccd1 vccd1 _7334_/D sky130_fd_sc_hd__nand3_1
X_6213_ _6213_/A _6213_/B vssd1 vssd1 vccd1 vccd1 _6215_/B sky130_fd_sc_hd__xnor2_1
X_4474_ _6599_/B vssd1 vssd1 vccd1 vccd1 _4723_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7193_ _7193_/A _7194_/B vssd1 vssd1 vccd1 vccd1 _7227_/A sky130_fd_sc_hd__nor2_1
X_6144_ _6142_/A _6128_/B _6128_/C vssd1 vssd1 vccd1 vccd1 _6145_/B sky130_fd_sc_hd__a21oi_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6075_ _6075_/A _6075_/B vssd1 vssd1 vccd1 vccd1 _6307_/B sky130_fd_sc_hd__nor2_1
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5026_ _5026_/A _5026_/B _5026_/C vssd1 vssd1 vccd1 vccd1 _5027_/B sky130_fd_sc_hd__and3_1
XFILLER_26_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6977_ _7199_/B _6947_/B _6977_/S vssd1 vssd1 vccd1 vccd1 _6978_/B sky130_fd_sc_hd__mux2_1
X_8716_ input3/X _8716_/D vssd1 vssd1 vccd1 vccd1 _8716_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5928_ _5949_/A _5949_/B vssd1 vssd1 vccd1 vccd1 _5929_/B sky130_fd_sc_hd__xor2_1
XFILLER_13_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8647_ input3/X _8647_/D vssd1 vssd1 vccd1 vccd1 _8647_/Q sky130_fd_sc_hd__dfxtp_1
X_5859_ _5859_/A _5859_/B vssd1 vssd1 vccd1 vccd1 _5862_/B sky130_fd_sc_hd__xor2_1
X_8578_ input3/X _8578_/D vssd1 vssd1 vccd1 vccd1 _8578_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7529_ _7529_/A _7537_/B vssd1 vssd1 vccd1 vccd1 _7532_/A sky130_fd_sc_hd__xnor2_1
XFILLER_79_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7880_ _7880_/A _7880_/B _7880_/C vssd1 vssd1 vccd1 vccd1 _7882_/B sky130_fd_sc_hd__nand3_1
X_6900_ _6900_/A vssd1 vssd1 vccd1 vccd1 _7135_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6831_ _7265_/A _6831_/B vssd1 vssd1 vccd1 vccd1 _6833_/A sky130_fd_sc_hd__nor2_1
XFILLER_50_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6762_ _7219_/A _7265_/A vssd1 vssd1 vccd1 vccd1 _6767_/A sky130_fd_sc_hd__nor2_1
X_8501_ _8501_/A _8501_/B vssd1 vssd1 vccd1 vccd1 _8502_/B sky130_fd_sc_hd__nand2_1
XFILLER_23_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6693_ _6670_/A _6673_/A _7249_/B vssd1 vssd1 vccd1 vccd1 _6703_/C sky130_fd_sc_hd__a21o_1
X_5713_ _5713_/A _5713_/B vssd1 vssd1 vccd1 vccd1 _5713_/Y sky130_fd_sc_hd__nand2_1
X_8432_ _8493_/A _8432_/B vssd1 vssd1 vccd1 vccd1 _8492_/A sky130_fd_sc_hd__nand2_1
X_5644_ _5953_/B _6042_/B vssd1 vssd1 vccd1 vccd1 _5701_/A sky130_fd_sc_hd__nor2_2
X_8363_ _8363_/A _8363_/B vssd1 vssd1 vccd1 vccd1 _8443_/B sky130_fd_sc_hd__xnor2_1
X_7314_ _7314_/A vssd1 vssd1 vccd1 vccd1 _7418_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_5575_ _5575_/A _6038_/A vssd1 vssd1 vccd1 vccd1 _5713_/A sky130_fd_sc_hd__nand2_1
X_8294_ _8294_/A _8294_/B vssd1 vssd1 vccd1 vccd1 _8295_/B sky130_fd_sc_hd__nand2_1
X_4526_ _5159_/A vssd1 vssd1 vccd1 vccd1 _4728_/B sky130_fd_sc_hd__clkbuf_2
X_4457_ _4459_/A vssd1 vssd1 vccd1 vccd1 _4457_/Y sky130_fd_sc_hd__inv_2
X_7245_ _7245_/A _7245_/B vssd1 vssd1 vccd1 vccd1 _7294_/A sky130_fd_sc_hd__nor2_1
XFILLER_104_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7176_ _7176_/A _7176_/B _7176_/C vssd1 vssd1 vccd1 vccd1 _7243_/A sky130_fd_sc_hd__and3_1
X_4388_ _4389_/A vssd1 vssd1 vccd1 vccd1 _4388_/Y sky130_fd_sc_hd__inv_2
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6127_ _6082_/B _5882_/A _6083_/C _6034_/B vssd1 vssd1 vccd1 vccd1 _6128_/C sky130_fd_sc_hd__o211a_1
XFILLER_100_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6058_ _6065_/A _6058_/B vssd1 vssd1 vccd1 vccd1 _6058_/X sky130_fd_sc_hd__and2_1
XFILLER_85_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5009_ _5132_/B _5009_/B vssd1 vssd1 vccd1 vccd1 _5014_/C sky130_fd_sc_hd__or2_1
XFILLER_45_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5360_ _8638_/Q _8637_/Q _5360_/C vssd1 vssd1 vccd1 vccd1 _5366_/C sky130_fd_sc_hd__and3_1
XFILLER_99_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5291_ _8619_/Q _5300_/B vssd1 vssd1 vccd1 vccd1 _5291_/X sky130_fd_sc_hd__or2_1
XFILLER_99_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7030_ _7417_/A _7030_/B vssd1 vssd1 vccd1 vccd1 _7032_/A sky130_fd_sc_hd__nand2_1
XFILLER_101_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7932_ _7929_/X _7930_/Y _7850_/X _7851_/Y vssd1 vssd1 vccd1 vccd1 _7938_/B sky130_fd_sc_hd__o211a_1
XFILLER_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7863_ _8209_/A _7764_/A _7877_/A vssd1 vssd1 vccd1 vccd1 _7865_/B sky130_fd_sc_hd__a21oi_1
XFILLER_70_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6814_ _6814_/A _6814_/B vssd1 vssd1 vccd1 vccd1 _6899_/A sky130_fd_sc_hd__xnor2_2
X_7794_ _8283_/A _7664_/X _7685_/X _7665_/A vssd1 vssd1 vccd1 vccd1 _7924_/B sky130_fd_sc_hd__a211o_1
XFILLER_50_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6745_ _6753_/B vssd1 vssd1 vccd1 vccd1 _6842_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_50_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8415_ _8415_/A _8415_/B _8415_/C vssd1 vssd1 vccd1 vccd1 _8416_/B sky130_fd_sc_hd__and3_1
X_6676_ _7249_/B _6700_/B _6769_/A _7296_/B _7418_/B vssd1 vssd1 vccd1 vccd1 _6676_/X
+ sky130_fd_sc_hd__a32o_1
X_5627_ _8652_/Q _7676_/A vssd1 vssd1 vccd1 vccd1 _5633_/B sky130_fd_sc_hd__and2b_1
X_8346_ _8346_/A _8355_/B vssd1 vssd1 vccd1 vccd1 _8347_/B sky130_fd_sc_hd__xnor2_1
X_5558_ _5558_/A _5724_/B _5794_/C vssd1 vssd1 vccd1 vccd1 _5595_/A sky130_fd_sc_hd__and3_1
X_8277_ _7817_/X _7816_/B _8445_/A _8245_/B _8276_/Y vssd1 vssd1 vccd1 vccd1 _8368_/B
+ sky130_fd_sc_hd__a41o_1
X_4509_ _8610_/Q vssd1 vssd1 vccd1 vccd1 _7676_/A sky130_fd_sc_hd__buf_4
X_7228_ _6773_/A _6862_/A _7222_/X vssd1 vssd1 vccd1 vccd1 _7229_/B sky130_fd_sc_hd__a21o_1
X_5489_ _5494_/A vssd1 vssd1 vccd1 vccd1 _5881_/B sky130_fd_sc_hd__clkbuf_2
X_7159_ _7159_/A _7159_/B vssd1 vssd1 vccd1 vccd1 _7212_/B sky130_fd_sc_hd__xnor2_1
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8785__63 vssd1 vssd1 vccd1 vccd1 _8785__63/HI _8894_/A sky130_fd_sc_hd__conb_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4860_ _4860_/A _4961_/B vssd1 vssd1 vccd1 vccd1 _5087_/A sky130_fd_sc_hd__nor2_1
X_4791_ _4848_/A _4795_/B vssd1 vssd1 vccd1 vccd1 _4872_/A sky130_fd_sc_hd__or2_1
XFILLER_32_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6530_ _6526_/A _6511_/X _6513_/X _6529_/Y vssd1 vssd1 vccd1 vccd1 _8691_/D sky130_fd_sc_hd__a22o_1
XFILLER_9_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6461_ _6463_/B _6461_/B _6461_/C vssd1 vssd1 vccd1 vccd1 _6462_/A sky130_fd_sc_hd__and3b_1
X_8200_ _8313_/A _8200_/B vssd1 vssd1 vccd1 vccd1 _8201_/B sky130_fd_sc_hd__nor2_1
X_5412_ _5412_/A vssd1 vssd1 vccd1 vccd1 _5412_/X sky130_fd_sc_hd__buf_2
X_6392_ _8683_/Q _6391_/X _8684_/Q vssd1 vssd1 vccd1 vccd1 _6393_/B sky130_fd_sc_hd__a21o_1
X_8131_ _8212_/B _8131_/B vssd1 vssd1 vccd1 vccd1 _8132_/B sky130_fd_sc_hd__nor2_1
X_5343_ _6475_/D _5342_/C _8633_/Q vssd1 vssd1 vccd1 vccd1 _5344_/B sky130_fd_sc_hd__a21o_1
XFILLER_99_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8062_ _7836_/B _8446_/S _8079_/B vssd1 vssd1 vccd1 vccd1 _8065_/A sky130_fd_sc_hd__o21ai_1
X_5274_ _8654_/Q _5271_/X _5272_/X _5273_/X vssd1 vssd1 vccd1 vccd1 _8612_/D sky130_fd_sc_hd__o211a_1
X_7013_ _7013_/A _7013_/B vssd1 vssd1 vccd1 vccd1 _7013_/Y sky130_fd_sc_hd__nand2_1
XFILLER_68_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7915_ _7920_/A _7985_/C vssd1 vssd1 vccd1 vccd1 _7984_/B sky130_fd_sc_hd__xnor2_1
XFILLER_55_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8895_ _8895_/A _4412_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[4] sky130_fd_sc_hd__ebufn_8
X_7846_ _8094_/A _7846_/B vssd1 vssd1 vccd1 vccd1 _7847_/A sky130_fd_sc_hd__and2_1
XFILLER_51_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7777_ _8395_/A _7853_/B _7777_/C vssd1 vssd1 vccd1 vccd1 _7850_/B sky130_fd_sc_hd__or3_1
X_4989_ _4989_/A vssd1 vssd1 vccd1 vccd1 _5143_/B sky130_fd_sc_hd__clkbuf_2
X_6728_ _6728_/A _7048_/B vssd1 vssd1 vccd1 vccd1 _6729_/B sky130_fd_sc_hd__nor2_1
XFILLER_11_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6659_ _6642_/X _6643_/X _6657_/A vssd1 vssd1 vccd1 vccd1 _7237_/C sky130_fd_sc_hd__a21oi_2
X_8329_ _8392_/A _8392_/B vssd1 vssd1 vccd1 vccd1 _8393_/B sky130_fd_sc_hd__xor2_1
XFILLER_11_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5961_ _5961_/A _5961_/B vssd1 vssd1 vccd1 vccd1 _5964_/B sky130_fd_sc_hd__or2_1
XFILLER_37_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7700_ _7699_/B _8546_/A vssd1 vssd1 vccd1 vccd1 _7701_/B sky130_fd_sc_hd__and2b_1
X_4912_ _5240_/B vssd1 vssd1 vccd1 vccd1 _5241_/A sky130_fd_sc_hd__clkbuf_2
X_8680_ input3/X _8680_/D vssd1 vssd1 vccd1 vccd1 _8680_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7631_ _8709_/Q _7631_/B vssd1 vssd1 vccd1 vccd1 _7631_/X sky130_fd_sc_hd__and2b_1
XFILLER_33_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5892_ _5507_/A _5506_/B _5507_/B _5549_/Y _5794_/A vssd1 vssd1 vccd1 vccd1 _5897_/B
+ sky130_fd_sc_hd__o311a_1
X_4843_ _4859_/A _4871_/A vssd1 vssd1 vccd1 vccd1 _5245_/C sky130_fd_sc_hd__nor2_1
XFILLER_20_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7562_ _8561_/A _8566_/A _7560_/X _7561_/X _4581_/A vssd1 vssd1 vccd1 vccd1 _8706_/D
+ sky130_fd_sc_hd__o311ai_1
XFILLER_20_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4774_ _5263_/A _4775_/C _4775_/A vssd1 vssd1 vccd1 vccd1 _4776_/B sky130_fd_sc_hd__a21o_1
X_7493_ _7493_/A _7509_/A vssd1 vssd1 vccd1 vccd1 _7493_/Y sky130_fd_sc_hd__nor2_1
X_6513_ _6513_/A vssd1 vssd1 vccd1 vccd1 _6513_/X sky130_fd_sc_hd__clkbuf_2
X_6444_ _6444_/A vssd1 vssd1 vccd1 vccd1 _8676_/D sky130_fd_sc_hd__clkbuf_1
X_6375_ _6375_/A _6375_/B vssd1 vssd1 vccd1 vccd1 _6375_/X sky130_fd_sc_hd__and2_1
X_8114_ _8317_/B _8027_/X _8026_/Y _8327_/A vssd1 vssd1 vccd1 vccd1 _8225_/A sky130_fd_sc_hd__a2bb2o_1
X_5326_ _8627_/Q _5324_/B _5325_/X vssd1 vssd1 vccd1 vccd1 _5327_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8045_ _8043_/Y _8044_/X _8031_/A vssd1 vssd1 vccd1 vccd1 _8158_/A sky130_fd_sc_hd__a21oi_2
X_5257_ _5070_/D _5087_/X _5252_/X _5256_/X vssd1 vssd1 vccd1 vccd1 _5257_/X sky130_fd_sc_hd__o31a_1
X_5188_ _5229_/D _5029_/B _5186_/X _5187_/X vssd1 vssd1 vccd1 vccd1 _5188_/X sky130_fd_sc_hd__o31a_1
XFILLER_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8755__33 vssd1 vssd1 vccd1 vccd1 _8755__33/HI _8850_/A sky130_fd_sc_hd__conb_1
X_8878_ _8878_/A _4397_/Y vssd1 vssd1 vccd1 vccd1 io_out[25] sky130_fd_sc_hd__ebufn_8
XFILLER_71_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7829_ _7829_/A _7829_/B vssd1 vssd1 vccd1 vccd1 _7830_/B sky130_fd_sc_hd__and2_1
XFILLER_51_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4490_ _4820_/A vssd1 vssd1 vccd1 vccd1 _4769_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6160_ _6163_/A _6164_/D vssd1 vssd1 vccd1 vccd1 _6311_/A sky130_fd_sc_hd__nand2_1
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5111_ _5111_/A _5111_/B vssd1 vssd1 vccd1 vccd1 _5111_/X sky130_fd_sc_hd__or2_1
XFILLER_85_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6091_ _6060_/A _6059_/B _6058_/X vssd1 vssd1 vccd1 vccd1 _6091_/X sky130_fd_sc_hd__o21ba_1
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5042_ _5042_/A _5193_/D vssd1 vssd1 vccd1 vccd1 _5046_/B sky130_fd_sc_hd__or2_1
XFILLER_53_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6993_ _6988_/X _6989_/Y _6853_/X _6894_/Y vssd1 vssd1 vccd1 vccd1 _6993_/Y sky130_fd_sc_hd__a211oi_2
XFILLER_53_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5944_ _5941_/A _5941_/B _5943_/Y vssd1 vssd1 vccd1 vccd1 _6170_/A sky130_fd_sc_hd__a21oi_1
XFILLER_80_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5875_ _5875_/A _5875_/B vssd1 vssd1 vccd1 vccd1 _5876_/B sky130_fd_sc_hd__xnor2_1
X_8663_ input3/X _8663_/D vssd1 vssd1 vccd1 vccd1 _8663_/Q sky130_fd_sc_hd__dfxtp_1
X_7614_ _7611_/A _7611_/C _7611_/B vssd1 vssd1 vccd1 vccd1 _7618_/A sky130_fd_sc_hd__a21bo_1
X_4826_ _4908_/A _4839_/B _4825_/Y _4864_/B vssd1 vssd1 vccd1 vccd1 _5119_/A sky130_fd_sc_hd__a2bb2o_1
X_8594_ input3/X _8594_/D vssd1 vssd1 vccd1 vccd1 _8594_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7545_ _7545_/A _7545_/B _7545_/C vssd1 vssd1 vccd1 vccd1 _7547_/B sky130_fd_sc_hd__or3_1
X_4757_ _8536_/A _4757_/B vssd1 vssd1 vccd1 vccd1 _4758_/A sky130_fd_sc_hd__and2_1
X_7476_ _7482_/A _7482_/B vssd1 vssd1 vccd1 vccd1 _7477_/B sky130_fd_sc_hd__or2_1
XFILLER_4_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4688_ _5259_/B _4707_/A vssd1 vssd1 vccd1 vccd1 _4688_/X sky130_fd_sc_hd__or2_1
X_6427_ _6468_/B vssd1 vssd1 vccd1 vccd1 _6427_/X sky130_fd_sc_hd__clkbuf_4
X_6358_ _6358_/A _6358_/B vssd1 vssd1 vccd1 vccd1 _6358_/X sky130_fd_sc_hd__or2_1
XFILLER_88_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5309_ _8641_/Q _8640_/Q _5309_/C vssd1 vssd1 vccd1 vccd1 _5309_/X sky130_fd_sc_hd__or3_1
XFILLER_102_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6289_ _6237_/A _6237_/B _6288_/X vssd1 vssd1 vccd1 vccd1 _6290_/B sky130_fd_sc_hd__a21oi_1
X_8028_ _7769_/A _8026_/Y _8027_/X vssd1 vssd1 vccd1 vccd1 _8029_/B sky130_fd_sc_hd__a21o_1
XFILLER_75_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5660_ _5660_/A vssd1 vssd1 vccd1 vccd1 _5660_/Y sky130_fd_sc_hd__inv_2
XFILLER_43_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4611_ _8578_/Q _4610_/C _8579_/Q vssd1 vssd1 vccd1 vccd1 _4612_/C sky130_fd_sc_hd__a21o_1
X_5591_ _5718_/A _5718_/B vssd1 vssd1 vccd1 vccd1 _5601_/A sky130_fd_sc_hd__xnor2_1
X_7330_ _7330_/A _7330_/B _7330_/C vssd1 vssd1 vccd1 vccd1 _7333_/A sky130_fd_sc_hd__and3_1
X_4542_ _4542_/A _4542_/B _4542_/C _4542_/D vssd1 vssd1 vccd1 vccd1 _4567_/B sky130_fd_sc_hd__and4_4
X_7261_ _7341_/A _7341_/B _7275_/B _7260_/B _7260_/A vssd1 vssd1 vccd1 vccd1 _7362_/A
+ sky130_fd_sc_hd__a32o_1
X_4473_ _7871_/A vssd1 vssd1 vccd1 vccd1 _6599_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_104_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6212_ _6008_/A _6008_/B _6013_/A vssd1 vssd1 vccd1 vccd1 _6249_/A sky130_fd_sc_hd__a21o_1
X_7192_ _7137_/B _6872_/B _6876_/A vssd1 vssd1 vccd1 vccd1 _7192_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_97_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6143_ _6323_/B _6143_/B vssd1 vssd1 vccd1 vccd1 _6322_/B sky130_fd_sc_hd__nor2_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6074_ _6074_/A _6074_/B _6074_/C vssd1 vssd1 vccd1 vccd1 _6075_/B sky130_fd_sc_hd__nor3_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5025_ _5180_/B vssd1 vssd1 vccd1 vccd1 _5151_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_72_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6976_ _7194_/B vssd1 vssd1 vccd1 vccd1 _7199_/B sky130_fd_sc_hd__inv_2
X_8715_ input3/X _8715_/D vssd1 vssd1 vccd1 vccd1 _8715_/Q sky130_fd_sc_hd__dfxtp_1
X_5927_ _5754_/B _5983_/A _5828_/B _5831_/A _5831_/B vssd1 vssd1 vccd1 vccd1 _5949_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_13_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5858_ _5858_/A _5858_/B vssd1 vssd1 vccd1 vccd1 _5859_/B sky130_fd_sc_hd__xor2_1
X_8646_ input3/X _8646_/D vssd1 vssd1 vccd1 vccd1 _8646_/Q sky130_fd_sc_hd__dfxtp_2
X_5789_ _5789_/A _5789_/B vssd1 vssd1 vccd1 vccd1 _5789_/Y sky130_fd_sc_hd__nand2_1
X_8577_ input3/X _8577_/D vssd1 vssd1 vccd1 vccd1 _8577_/Q sky130_fd_sc_hd__dfxtp_1
X_4809_ _5092_/C _5241_/C vssd1 vssd1 vccd1 vccd1 _5009_/B sky130_fd_sc_hd__or2_1
XFILLER_21_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7528_ _6711_/A _5325_/X _6513_/A _7527_/X vssd1 vssd1 vccd1 vccd1 _8702_/D sky130_fd_sc_hd__a22o_1
XFILLER_5_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7459_ _7459_/A _7459_/B vssd1 vssd1 vccd1 vccd1 _7485_/B sky130_fd_sc_hd__nor2_1
XFILLER_79_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6830_ _6767_/A _6767_/B _6829_/X vssd1 vssd1 vccd1 vccd1 _6834_/A sky130_fd_sc_hd__a21oi_1
XFILLER_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6761_ _7179_/A vssd1 vssd1 vccd1 vccd1 _7265_/A sky130_fd_sc_hd__clkbuf_2
X_8500_ _8500_/A _8500_/B _8500_/C vssd1 vssd1 vccd1 vccd1 _8501_/B sky130_fd_sc_hd__or3_1
X_5712_ _5783_/A _5712_/B vssd1 vssd1 vccd1 vccd1 _6061_/B sky130_fd_sc_hd__nor2_1
X_6692_ _6692_/A _6692_/B vssd1 vssd1 vccd1 vccd1 _6705_/A sky130_fd_sc_hd__xnor2_2
XFILLER_31_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8431_ _8431_/A _8431_/B vssd1 vssd1 vccd1 vccd1 _8432_/B sky130_fd_sc_hd__or2_1
X_5643_ _5643_/A _5643_/B vssd1 vssd1 vccd1 vccd1 _6042_/B sky130_fd_sc_hd__xor2_4
X_8362_ _8361_/Y _8304_/B _8302_/X vssd1 vssd1 vccd1 vccd1 _8364_/A sky130_fd_sc_hd__a21boi_1
X_5574_ _6082_/B _5574_/B _5575_/A _5574_/D vssd1 vssd1 vccd1 vccd1 _6038_/A sky130_fd_sc_hd__nand4_1
X_7313_ _7313_/A _7313_/B vssd1 vssd1 vccd1 vccd1 _7325_/A sky130_fd_sc_hd__xnor2_1
X_4525_ _5185_/A vssd1 vssd1 vccd1 vccd1 _5159_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_8293_ _8293_/A _8248_/B vssd1 vssd1 vccd1 vccd1 _8294_/B sky130_fd_sc_hd__or2b_1
X_7244_ _7315_/A _7299_/B vssd1 vssd1 vccd1 vccd1 _7248_/B sky130_fd_sc_hd__xnor2_1
X_4456_ _4456_/A vssd1 vssd1 vccd1 vccd1 _4456_/Y sky130_fd_sc_hd__inv_2
X_4387_ _4389_/A vssd1 vssd1 vccd1 vccd1 _4387_/Y sky130_fd_sc_hd__inv_2
X_7175_ _7175_/A _7175_/B vssd1 vssd1 vccd1 vccd1 _7315_/A sky130_fd_sc_hd__nor2_2
X_6126_ _5954_/A _6111_/S _5964_/B _6124_/Y _6125_/X vssd1 vssd1 vccd1 vccd1 _6128_/B
+ sky130_fd_sc_hd__a32o_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6057_ _6057_/A _6057_/B vssd1 vssd1 vccd1 vccd1 _6058_/B sky130_fd_sc_hd__nand2_1
XFILLER_66_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5008_ _5185_/C _5029_/B _5180_/B vssd1 vssd1 vccd1 vccd1 _5047_/B sky130_fd_sc_hd__or3_1
XFILLER_14_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6959_ _7010_/A _7004_/C vssd1 vssd1 vccd1 vccd1 _6960_/B sky130_fd_sc_hd__nand2_1
XFILLER_53_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8629_ input3/X _8629_/D vssd1 vssd1 vccd1 vccd1 _8629_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5290_ _5290_/A vssd1 vssd1 vccd1 vccd1 _5300_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_4_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7931_ _7850_/X _7851_/Y _7929_/X _7930_/Y vssd1 vssd1 vccd1 vccd1 _7938_/A sky130_fd_sc_hd__a211oi_2
XFILLER_27_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7862_ _7862_/A _7862_/B vssd1 vssd1 vccd1 vccd1 _7877_/A sky130_fd_sc_hd__nor2_2
XFILLER_51_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6813_ _7048_/A _7046_/A vssd1 vssd1 vccd1 vccd1 _6814_/B sky130_fd_sc_hd__nor2_1
X_7793_ _7902_/A _7902_/B vssd1 vssd1 vccd1 vccd1 _7924_/A sky130_fd_sc_hd__xnor2_1
XFILLER_35_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6744_ _6744_/A _6772_/A vssd1 vssd1 vccd1 vccd1 _6753_/B sky130_fd_sc_hd__nand2_2
X_6675_ _6697_/B vssd1 vssd1 vccd1 vccd1 _7296_/B sky130_fd_sc_hd__clkbuf_2
X_8414_ _8415_/A _8415_/B _8415_/C vssd1 vssd1 vccd1 vccd1 _8416_/A sky130_fd_sc_hd__a21oi_1
X_5626_ _5679_/A _5680_/A _5680_/B _5624_/X _5641_/A vssd1 vssd1 vccd1 vccd1 _5631_/B
+ sky130_fd_sc_hd__a311o_1
X_8345_ _8376_/A _8345_/B vssd1 vssd1 vccd1 vccd1 _8355_/B sky130_fd_sc_hd__xnor2_1
X_5557_ _5577_/B _5556_/C _5556_/A vssd1 vssd1 vccd1 vccd1 _5569_/B sky130_fd_sc_hd__a21oi_1
XFILLER_104_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8276_ _8437_/A _8276_/B vssd1 vssd1 vccd1 vccd1 _8276_/Y sky130_fd_sc_hd__nor2_1
X_4508_ _4850_/A _4822_/A _4507_/X vssd1 vssd1 vccd1 vccd1 _4518_/C sky130_fd_sc_hd__o21a_1
X_5488_ _5539_/A _5533_/B vssd1 vssd1 vccd1 vccd1 _5488_/Y sky130_fd_sc_hd__nand2_1
X_4439_ _4451_/A vssd1 vssd1 vccd1 vccd1 _4444_/A sky130_fd_sc_hd__clkbuf_2
X_7227_ _7227_/A _7425_/B vssd1 vssd1 vccd1 vccd1 _7231_/A sky130_fd_sc_hd__nand2_1
X_7158_ _7158_/A _7158_/B vssd1 vssd1 vccd1 vccd1 _7469_/A sky130_fd_sc_hd__xnor2_4
XFILLER_86_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7089_ _7456_/A vssd1 vssd1 vccd1 vccd1 _7462_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_100_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6109_ _6109_/A _6109_/B vssd1 vssd1 vccd1 vccd1 _6125_/A sky130_fd_sc_hd__nor2_1
XFILLER_27_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4790_ _7631_/B _4822_/C vssd1 vssd1 vccd1 vccd1 _4795_/B sky130_fd_sc_hd__and2_1
XFILLER_60_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6460_ _8680_/Q _6459_/B _6454_/B _8682_/Q vssd1 vssd1 vccd1 vccd1 _6461_/C sky130_fd_sc_hd__a31o_1
X_5411_ _5411_/A vssd1 vssd1 vccd1 vccd1 _8647_/D sky130_fd_sc_hd__clkbuf_1
X_6391_ _8680_/Q _6459_/B _6398_/A _6390_/X _8682_/Q vssd1 vssd1 vccd1 vccd1 _6391_/X
+ sky130_fd_sc_hd__a221o_1
X_8130_ _8225_/A _8130_/B vssd1 vssd1 vccd1 vccd1 _8131_/B sky130_fd_sc_hd__nor2_1
X_5342_ _8633_/Q _8632_/Q _5342_/C vssd1 vssd1 vccd1 vccd1 _5346_/B sky130_fd_sc_hd__and3_1
X_8061_ _7790_/A _8166_/A _8296_/A vssd1 vssd1 vccd1 vccd1 _8079_/B sky130_fd_sc_hd__a21o_1
XFILLER_99_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7012_ _7012_/A _7012_/B vssd1 vssd1 vccd1 vccd1 _7149_/B sky130_fd_sc_hd__xor2_2
X_5273_ _5296_/A vssd1 vssd1 vccd1 vccd1 _5273_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_99_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7914_ _8296_/A _7911_/Y _8006_/A vssd1 vssd1 vccd1 vccd1 _7985_/C sky130_fd_sc_hd__a21oi_2
X_8894_ _8894_/A _4414_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[3] sky130_fd_sc_hd__ebufn_8
X_7845_ _7845_/A _7849_/A vssd1 vssd1 vccd1 vccd1 _7846_/B sky130_fd_sc_hd__nand2_1
XFILLER_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7776_ _7862_/A vssd1 vssd1 vccd1 vccd1 _8395_/A sky130_fd_sc_hd__buf_2
X_4988_ _4988_/A _5074_/B vssd1 vssd1 vccd1 vccd1 _5219_/D sky130_fd_sc_hd__or2_2
X_6727_ _7245_/B vssd1 vssd1 vccd1 vccd1 _7048_/B sky130_fd_sc_hd__clkbuf_2
X_6658_ _7237_/B vssd1 vssd1 vccd1 vccd1 _6798_/B sky130_fd_sc_hd__clkbuf_2
X_5609_ _6042_/A vssd1 vssd1 vccd1 vccd1 _6323_/C sky130_fd_sc_hd__buf_2
X_8328_ _8331_/B _8328_/B vssd1 vssd1 vccd1 vccd1 _8392_/B sky130_fd_sc_hd__xor2_1
X_6589_ _6744_/A _7425_/A _6588_/C vssd1 vssd1 vccd1 vccd1 _6589_/X sky130_fd_sc_hd__a21o_1
XFILLER_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8259_ _8269_/A _8269_/B vssd1 vssd1 vccd1 vccd1 _8260_/B sky130_fd_sc_hd__xor2_1
XFILLER_59_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5960_ _5870_/B _5986_/A _5968_/B _5983_/B vssd1 vssd1 vccd1 vccd1 _6178_/A sky130_fd_sc_hd__a22o_1
XFILLER_52_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4911_ _4975_/B _5114_/B vssd1 vssd1 vccd1 vccd1 _5240_/B sky130_fd_sc_hd__nand2_2
X_5891_ _5889_/X _5814_/B _5890_/X vssd1 vssd1 vccd1 vccd1 _5915_/A sky130_fd_sc_hd__o21bai_1
X_7630_ _8709_/Q _8606_/Q vssd1 vssd1 vccd1 vccd1 _7654_/B sky130_fd_sc_hd__xnor2_4
X_4842_ _4849_/A _4850_/B _4842_/C _4824_/B vssd1 vssd1 vccd1 vccd1 _4871_/A sky130_fd_sc_hd__or4b_2
XFILLER_20_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7561_ _7875_/A _7552_/A _8552_/B vssd1 vssd1 vccd1 vccd1 _7561_/X sky130_fd_sc_hd__a21o_1
X_4773_ _4773_/A vssd1 vssd1 vccd1 vccd1 _8608_/D sky130_fd_sc_hd__clkbuf_1
X_7492_ _7492_/A _7492_/B _7492_/C _7492_/D vssd1 vssd1 vccd1 vccd1 _7509_/A sky130_fd_sc_hd__or4_2
X_6512_ _6512_/A vssd1 vssd1 vccd1 vccd1 _6513_/A sky130_fd_sc_hd__clkbuf_2
X_6443_ _6445_/B _6443_/B _6461_/B vssd1 vssd1 vccd1 vccd1 _6444_/A sky130_fd_sc_hd__and3b_1
X_6374_ _5413_/X _6373_/Y _6371_/A _4582_/B vssd1 vssd1 vccd1 vccd1 _8663_/D sky130_fd_sc_hd__o2bb2a_1
X_8113_ _8205_/B _8113_/B vssd1 vssd1 vccd1 vccd1 _8120_/A sky130_fd_sc_hd__xnor2_2
X_5325_ _6511_/A vssd1 vssd1 vccd1 vccd1 _5325_/X sky130_fd_sc_hd__buf_2
X_8044_ _8044_/A _7975_/B vssd1 vssd1 vccd1 vccd1 _8044_/X sky130_fd_sc_hd__or2b_1
X_5256_ _5256_/A _5256_/B _5256_/C _5256_/D vssd1 vssd1 vccd1 vccd1 _5256_/X sky130_fd_sc_hd__or4_1
X_5187_ _4885_/X _5132_/B _5180_/X _5027_/B _4731_/A vssd1 vssd1 vccd1 vccd1 _5187_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_56_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8877_ _8877_/A _4395_/Y vssd1 vssd1 vccd1 vccd1 io_out[24] sky130_fd_sc_hd__ebufn_8
XFILLER_36_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7828_ _7829_/A _7829_/B vssd1 vssd1 vccd1 vccd1 _7830_/A sky130_fd_sc_hd__nor2_1
XFILLER_24_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8770__48 vssd1 vssd1 vccd1 vccd1 _8770__48/HI _8879_/A sky130_fd_sc_hd__conb_1
X_7759_ _7759_/A _7759_/B vssd1 vssd1 vccd1 vccd1 _7853_/C sky130_fd_sc_hd__xor2_1
XFILLER_7_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5110_ _5241_/A _5110_/B _5202_/B _5110_/D vssd1 vssd1 vccd1 vccd1 _5111_/B sky130_fd_sc_hd__or4_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6090_ _6135_/A vssd1 vssd1 vccd1 vccd1 _6090_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5041_ _5041_/A _5041_/B vssd1 vssd1 vccd1 vccd1 _5245_/D sky130_fd_sc_hd__nor2_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6992_ _6992_/A _6893_/A vssd1 vssd1 vccd1 vccd1 _6992_/X sky130_fd_sc_hd__or2b_1
X_5943_ _5943_/A _5943_/B vssd1 vssd1 vccd1 vccd1 _5943_/Y sky130_fd_sc_hd__nor2_1
X_5874_ _5991_/A _5874_/B vssd1 vssd1 vccd1 vccd1 _5875_/B sky130_fd_sc_hd__or2_1
X_8662_ input3/X _8662_/D vssd1 vssd1 vccd1 vccd1 _8662_/Q sky130_fd_sc_hd__dfxtp_1
X_7613_ _8712_/Q _6427_/X _7612_/X vssd1 vssd1 vccd1 vccd1 _8712_/D sky130_fd_sc_hd__a21bo_1
X_4825_ _4836_/B vssd1 vssd1 vccd1 vccd1 _4825_/Y sky130_fd_sc_hd__inv_2
X_8593_ input3/X _8593_/D vssd1 vssd1 vccd1 vccd1 _8593_/Q sky130_fd_sc_hd__dfxtp_1
X_7544_ _7529_/A _7532_/B _7538_/B _7543_/X vssd1 vssd1 vccd1 vccd1 _7545_/C sky130_fd_sc_hd__o31a_1
X_4756_ _4675_/B _4856_/A _4754_/X _5290_/A _4507_/X vssd1 vssd1 vccd1 vccd1 _4757_/B
+ sky130_fd_sc_hd__a32o_1
X_7475_ _7508_/A _7505_/B _7474_/X vssd1 vssd1 vccd1 vccd1 _7492_/B sky130_fd_sc_hd__o21a_1
X_4687_ _5259_/B _4707_/A vssd1 vssd1 vccd1 vccd1 _4695_/A sky130_fd_sc_hd__nand2_1
X_6426_ _6430_/A _6430_/C vssd1 vssd1 vccd1 vccd1 _6429_/A sky130_fd_sc_hd__and2_1
X_6357_ _6357_/A _6364_/B vssd1 vssd1 vccd1 vccd1 _6358_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5308_ _8637_/Q _5307_/X _8639_/Q _8638_/Q vssd1 vssd1 vccd1 vccd1 _5309_/C sky130_fd_sc_hd__o211a_1
XFILLER_0_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6288_ _6236_/B _6288_/B vssd1 vssd1 vccd1 vccd1 _6288_/X sky130_fd_sc_hd__and2b_1
XFILLER_102_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8027_ _8125_/A _7957_/C _7957_/D _8115_/A _7884_/A vssd1 vssd1 vccd1 vccd1 _8027_/X
+ sky130_fd_sc_hd__o32a_1
X_5239_ _5253_/B _5239_/B vssd1 vssd1 vccd1 vccd1 _5248_/B sky130_fd_sc_hd__or2_1
XFILLER_102_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8815__93 vssd1 vssd1 vccd1 vccd1 _8815__93/HI _8924_/A sky130_fd_sc_hd__conb_1
XFILLER_68_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4610_ _8578_/Q _8579_/Q _4610_/C vssd1 vssd1 vccd1 vccd1 _4614_/B sky130_fd_sc_hd__and3_1
X_5590_ _5590_/A _5590_/B vssd1 vssd1 vccd1 vccd1 _5718_/B sky130_fd_sc_hd__xnor2_1
X_4541_ _4789_/A _4541_/B _4541_/C _4861_/A vssd1 vssd1 vccd1 vccd1 _4542_/D sky130_fd_sc_hd__or4_1
X_7260_ _7260_/A _7260_/B vssd1 vssd1 vccd1 vccd1 _7275_/B sky130_fd_sc_hd__xor2_1
X_4472_ _8601_/Q vssd1 vssd1 vccd1 vccd1 _7871_/A sky130_fd_sc_hd__clkbuf_4
X_7191_ _7191_/A _7208_/A vssd1 vssd1 vccd1 vccd1 _7278_/A sky130_fd_sc_hd__xnor2_1
X_6211_ _6021_/A _6021_/B _6210_/X vssd1 vssd1 vccd1 vccd1 _6288_/B sky130_fd_sc_hd__a21bo_1
X_6142_ _6142_/A _6142_/B vssd1 vssd1 vccd1 vccd1 _6302_/A sky130_fd_sc_hd__xor2_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6073_ _6103_/A _6103_/B _6103_/C vssd1 vssd1 vccd1 vccd1 _6167_/A sky130_fd_sc_hd__o21ai_2
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5024_ _5118_/B _5182_/C _4916_/B _5183_/S vssd1 vssd1 vccd1 vccd1 _5024_/X sky130_fd_sc_hd__o31a_1
XFILLER_93_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6975_ _7107_/A _6881_/Y _6884_/B _6978_/A vssd1 vssd1 vccd1 vccd1 _6980_/A sky130_fd_sc_hd__a22o_1
XFILLER_80_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8714_ input3/X _8714_/D vssd1 vssd1 vccd1 vccd1 _8714_/Q sky130_fd_sc_hd__dfxtp_1
X_5926_ _6270_/A _5926_/B vssd1 vssd1 vccd1 vccd1 _5949_/A sky130_fd_sc_hd__xnor2_1
XFILLER_13_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8645_ input3/X _8645_/D vssd1 vssd1 vccd1 vccd1 _8645_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5857_ _5857_/A _5857_/B vssd1 vssd1 vccd1 vccd1 _5858_/B sky130_fd_sc_hd__nand2_1
X_8740__18 vssd1 vssd1 vccd1 vccd1 _8740__18/HI _8835_/A sky130_fd_sc_hd__conb_1
X_5788_ _5744_/A _5744_/B _5739_/A _5739_/B vssd1 vssd1 vccd1 vccd1 _5867_/A sky130_fd_sc_hd__o2bb2a_1
X_4808_ _4899_/A vssd1 vssd1 vccd1 vccd1 _5241_/C sky130_fd_sc_hd__clkbuf_2
X_8576_ input3/X _8576_/D vssd1 vssd1 vccd1 vccd1 _8576_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7527_ _7527_/A _7527_/B vssd1 vssd1 vccd1 vccd1 _7527_/X sky130_fd_sc_hd__xor2_1
X_4739_ _4739_/A _4739_/B vssd1 vssd1 vccd1 vccd1 _4760_/A sky130_fd_sc_hd__and2_1
X_7458_ _7458_/A _7458_/B _7458_/C vssd1 vssd1 vccd1 vccd1 _7459_/B sky130_fd_sc_hd__and3_1
X_6409_ _6400_/A _6409_/B _6409_/C vssd1 vssd1 vccd1 vccd1 _6410_/A sky130_fd_sc_hd__and3b_1
X_7389_ _7388_/A _7409_/A vssd1 vssd1 vccd1 vccd1 _7393_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6760_ _6760_/A _6705_/A vssd1 vssd1 vccd1 vccd1 _6878_/A sky130_fd_sc_hd__or2b_1
XFILLER_35_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5711_ _5861_/A _5711_/B _5711_/C vssd1 vssd1 vccd1 vccd1 _5712_/B sky130_fd_sc_hd__and3_1
X_6691_ _6719_/A _6691_/B vssd1 vssd1 vccd1 vccd1 _6692_/B sky130_fd_sc_hd__xnor2_2
X_8430_ _8431_/A _8431_/B vssd1 vssd1 vccd1 vccd1 _8493_/A sky130_fd_sc_hd__nand2_1
X_5642_ _5642_/A _5642_/B vssd1 vssd1 vccd1 vccd1 _5643_/B sky130_fd_sc_hd__nand2_2
X_8361_ _8361_/A vssd1 vssd1 vccd1 vccd1 _8361_/Y sky130_fd_sc_hd__inv_2
X_5573_ _5576_/B _5571_/C _5571_/A vssd1 vssd1 vccd1 vccd1 _5574_/D sky130_fd_sc_hd__a21o_1
X_7312_ _7332_/A _7332_/B _7311_/X vssd1 vssd1 vccd1 vccd1 _7390_/A sky130_fd_sc_hd__a21oi_1
X_4524_ _8594_/Q vssd1 vssd1 vccd1 vccd1 _5185_/A sky130_fd_sc_hd__clkbuf_2
X_8292_ _8292_/A _8292_/B vssd1 vssd1 vccd1 vccd1 _8294_/A sky130_fd_sc_hd__nand2_1
X_4455_ _4456_/A vssd1 vssd1 vccd1 vccd1 _4455_/Y sky130_fd_sc_hd__inv_2
X_7243_ _7243_/A vssd1 vssd1 vccd1 vccd1 _7296_/C sky130_fd_sc_hd__clkbuf_2
X_4386_ _4389_/A vssd1 vssd1 vccd1 vccd1 _4386_/Y sky130_fd_sc_hd__inv_2
X_7174_ _7417_/A _7174_/B vssd1 vssd1 vccd1 vccd1 _7254_/A sky130_fd_sc_hd__nor2_1
XFILLER_100_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6125_ _6125_/A _6125_/B vssd1 vssd1 vccd1 vccd1 _6125_/X sky130_fd_sc_hd__or2_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6056_ _6057_/A _6057_/B vssd1 vssd1 vccd1 vccd1 _6065_/A sky130_fd_sc_hd__or2_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5007_ _5007_/A vssd1 vssd1 vccd1 vccd1 _5029_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_38_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6958_ _7088_/A _7139_/A vssd1 vssd1 vccd1 vccd1 _7004_/C sky130_fd_sc_hd__nand2_1
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6889_ _6868_/A _6868_/B _6888_/X vssd1 vssd1 vccd1 vccd1 _6890_/B sky130_fd_sc_hd__o21a_1
XFILLER_22_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5909_ _5909_/A _6229_/A vssd1 vssd1 vccd1 vccd1 _5910_/B sky130_fd_sc_hd__or2_1
X_8628_ input3/X _8628_/D vssd1 vssd1 vccd1 vccd1 _8628_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8559_ _8566_/A _8552_/B _8567_/S vssd1 vssd1 vccd1 vccd1 _8563_/A sky130_fd_sc_hd__a21o_1
XFILLER_30_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7930_ _7929_/A _7929_/B _7929_/C vssd1 vssd1 vccd1 vccd1 _7930_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_82_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7861_ _8134_/A _7957_/C _7957_/D vssd1 vssd1 vccd1 vccd1 _7889_/A sky130_fd_sc_hd__or3_1
X_6812_ _6950_/A _6812_/B vssd1 vssd1 vccd1 vccd1 _6819_/A sky130_fd_sc_hd__xnor2_1
XFILLER_35_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7792_ _7796_/B _7792_/B vssd1 vssd1 vccd1 vccd1 _7902_/B sky130_fd_sc_hd__xnor2_1
XFILLER_51_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6743_ _7174_/B vssd1 vssd1 vccd1 vccd1 _7236_/B sky130_fd_sc_hd__buf_2
X_6674_ _6674_/A _6674_/B vssd1 vssd1 vccd1 vccd1 _6697_/B sky130_fd_sc_hd__xnor2_1
XFILLER_31_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8413_ _8412_/A _8409_/X _8471_/A _8412_/Y vssd1 vssd1 vccd1 vccd1 _8415_/C sky130_fd_sc_hd__a2bb2o_1
X_5625_ _8651_/Q _8609_/Q vssd1 vssd1 vccd1 vccd1 _5641_/A sky130_fd_sc_hd__and2b_1
X_8344_ _8377_/A _8377_/B vssd1 vssd1 vccd1 vccd1 _8345_/B sky130_fd_sc_hd__xor2_1
X_5556_ _5556_/A _5577_/B _5556_/C vssd1 vssd1 vccd1 vccd1 _5569_/A sky130_fd_sc_hd__and3_1
X_8275_ _8301_/B vssd1 vssd1 vccd1 vccd1 _8445_/A sky130_fd_sc_hd__clkbuf_2
X_4507_ _4849_/A vssd1 vssd1 vccd1 vccd1 _4507_/X sky130_fd_sc_hd__clkbuf_2
X_5487_ _5539_/A vssd1 vssd1 vccd1 vccd1 _6213_/A sky130_fd_sc_hd__buf_2
XFILLER_104_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4438_ _4438_/A vssd1 vssd1 vccd1 vccd1 _4438_/Y sky130_fd_sc_hd__inv_2
X_7226_ _7226_/A _7226_/B vssd1 vssd1 vccd1 vccd1 _7425_/B sky130_fd_sc_hd__nor2_1
XFILLER_104_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7157_ _7157_/A _7157_/B vssd1 vssd1 vccd1 vccd1 _7158_/B sky130_fd_sc_hd__xnor2_4
X_4369_ _4370_/A vssd1 vssd1 vccd1 vccd1 _4369_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7088_ _7088_/A _7088_/B vssd1 vssd1 vccd1 vccd1 _7456_/A sky130_fd_sc_hd__nand2_2
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6108_ _6108_/A vssd1 vssd1 vccd1 vccd1 _6109_/A sky130_fd_sc_hd__inv_2
XFILLER_46_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6039_ _6038_/A _6038_/C _6038_/B vssd1 vssd1 vccd1 vccd1 _6059_/B sky130_fd_sc_hd__a21oi_1
XFILLER_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8776__54 vssd1 vssd1 vccd1 vccd1 _8776__54/HI _8885_/A sky130_fd_sc_hd__conb_1
XFILLER_17_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5410_ _5412_/A _5413_/A _5607_/A vssd1 vssd1 vccd1 vccd1 _5411_/A sky130_fd_sc_hd__mux2_1
X_6390_ _8677_/Q _6388_/X _6450_/B vssd1 vssd1 vccd1 vccd1 _6390_/X sky130_fd_sc_hd__a21o_1
X_5341_ _6475_/D _5342_/C _5340_/Y vssd1 vssd1 vccd1 vccd1 _8632_/D sky130_fd_sc_hd__a21oi_1
X_8060_ _8060_/A _8060_/B vssd1 vssd1 vccd1 vccd1 _8446_/S sky130_fd_sc_hd__nand2_2
XFILLER_99_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7011_ _7011_/A _7011_/B vssd1 vssd1 vccd1 vccd1 _7012_/B sky130_fd_sc_hd__nand2_1
X_5272_ _8612_/Q _5275_/B vssd1 vssd1 vccd1 vccd1 _5272_/X sky130_fd_sc_hd__or2_1
XFILLER_95_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7913_ _7786_/A _7786_/B _8455_/A vssd1 vssd1 vccd1 vccd1 _8006_/A sky130_fd_sc_hd__o21ba_2
XFILLER_83_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8893_ _8893_/A _4417_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[2] sky130_fd_sc_hd__ebufn_8
XFILLER_70_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7844_ _7845_/A _7849_/A vssd1 vssd1 vccd1 vccd1 _8094_/A sky130_fd_sc_hd__or2_1
XFILLER_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7775_ _7775_/A _7852_/B vssd1 vssd1 vccd1 vccd1 _7850_/A sky130_fd_sc_hd__xor2_1
XFILLER_51_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6726_ _7249_/B vssd1 vssd1 vccd1 vccd1 _6728_/A sky130_fd_sc_hd__clkbuf_2
X_4987_ _5219_/A _5167_/B _4987_/C _4987_/D vssd1 vssd1 vccd1 vccd1 _4987_/X sky130_fd_sc_hd__or4_1
X_6657_ _6657_/A _6657_/B _6657_/C vssd1 vssd1 vccd1 vccd1 _7237_/B sky130_fd_sc_hd__and3_1
X_6588_ _6744_/A _7425_/A _6588_/C vssd1 vssd1 vccd1 vccd1 _6590_/A sky130_fd_sc_hd__and3_1
X_5608_ _5657_/A _5645_/B vssd1 vssd1 vccd1 vccd1 _6042_/A sky130_fd_sc_hd__and2_1
X_8327_ _8327_/A _8334_/A vssd1 vssd1 vccd1 vccd1 _8328_/B sky130_fd_sc_hd__xor2_1
X_5539_ _5539_/A _5539_/B _5580_/B vssd1 vssd1 vccd1 vccd1 _5578_/A sky130_fd_sc_hd__or3_1
X_8258_ _8258_/A _8258_/B vssd1 vssd1 vccd1 vccd1 _8269_/B sky130_fd_sc_hd__xnor2_1
XFILLER_78_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7209_ _7278_/A _7278_/B _7208_/X vssd1 vssd1 vccd1 vccd1 _7212_/A sky130_fd_sc_hd__a21bo_1
X_8189_ _8189_/A _8164_/B vssd1 vssd1 vccd1 vccd1 _8189_/X sky130_fd_sc_hd__or2b_1
XFILLER_86_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4910_ _5011_/A _5010_/B vssd1 vssd1 vccd1 vccd1 _5114_/B sky130_fd_sc_hd__or2_1
X_5890_ _5889_/B _5890_/B vssd1 vssd1 vccd1 vccd1 _5890_/X sky130_fd_sc_hd__and2b_1
X_4841_ _5094_/A _5101_/A vssd1 vssd1 vccd1 vccd1 _4933_/A sky130_fd_sc_hd__or2_1
X_7560_ _7875_/A _7552_/Y _7556_/X _7559_/X vssd1 vssd1 vccd1 vccd1 _7560_/X sky130_fd_sc_hd__o31a_1
X_4772_ _7547_/A _4772_/B _4772_/C vssd1 vssd1 vccd1 vccd1 _4773_/A sky130_fd_sc_hd__and3_1
X_7491_ _7487_/X _7488_/B _7489_/X _7490_/Y vssd1 vssd1 vccd1 vccd1 _7492_/D sky130_fd_sc_hd__a22o_1
X_6511_ _6511_/A vssd1 vssd1 vccd1 vccd1 _6511_/X sky130_fd_sc_hd__clkbuf_2
X_6442_ _6441_/B _8674_/Q _6435_/A _8676_/Q vssd1 vssd1 vccd1 vccd1 _6443_/B sky130_fd_sc_hd__a31o_1
X_8112_ _8134_/B _8126_/B vssd1 vssd1 vccd1 vccd1 _8113_/B sky130_fd_sc_hd__xnor2_2
X_6373_ _6373_/A _6373_/B vssd1 vssd1 vccd1 vccd1 _6373_/Y sky130_fd_sc_hd__xnor2_1
X_5324_ _8627_/Q _5324_/B vssd1 vssd1 vccd1 vccd1 _5330_/C sky130_fd_sc_hd__and2_1
XFILLER_102_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8043_ _8043_/A _8043_/B vssd1 vssd1 vccd1 vccd1 _8043_/Y sky130_fd_sc_hd__nand2_1
X_5255_ _5119_/A _5104_/B _5105_/A vssd1 vssd1 vccd1 vccd1 _5256_/D sky130_fd_sc_hd__o21a_1
XFILLER_57_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5186_ _4990_/A _5153_/A _5182_/C _5135_/C _4941_/C vssd1 vssd1 vccd1 vccd1 _5186_/X
+ sky130_fd_sc_hd__o41a_1
XFILLER_83_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8876_ _8876_/A _4394_/Y vssd1 vssd1 vccd1 vccd1 io_out[23] sky130_fd_sc_hd__ebufn_8
XFILLER_71_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7827_ _8134_/A _7777_/C _7841_/A _7841_/B vssd1 vssd1 vccd1 vccd1 _7829_/B sky130_fd_sc_hd__o22a_1
XFILLER_24_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7758_ _7758_/A _7886_/C vssd1 vssd1 vccd1 vccd1 _7759_/B sky130_fd_sc_hd__xnor2_1
X_6709_ _6765_/B _6709_/B vssd1 vssd1 vccd1 vccd1 _6789_/A sky130_fd_sc_hd__nand2_1
X_7689_ _8723_/Q _7689_/B vssd1 vssd1 vccd1 vccd1 _7690_/B sky130_fd_sc_hd__and2_1
XFILLER_7_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8746__24 vssd1 vssd1 vccd1 vccd1 _8746__24/HI _8841_/A sky130_fd_sc_hd__conb_1
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5040_ _5040_/A _5137_/B _5040_/C _4940_/Y vssd1 vssd1 vccd1 vccd1 _5040_/X sky130_fd_sc_hd__or4b_1
XFILLER_84_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6991_ _6991_/A _6892_/A vssd1 vssd1 vccd1 vccd1 _6991_/X sky130_fd_sc_hd__or2b_1
XFILLER_38_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5942_ _6074_/A _6074_/B _6074_/C vssd1 vssd1 vccd1 vccd1 _6075_/A sky130_fd_sc_hd__o21a_1
X_5873_ _6205_/A _5873_/B vssd1 vssd1 vccd1 vccd1 _5874_/B sky130_fd_sc_hd__nor2_1
X_8661_ input3/X _8661_/D vssd1 vssd1 vccd1 vccd1 _8661_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7612_ _8557_/A _8568_/A _7612_/C _7622_/S vssd1 vssd1 vccd1 vccd1 _7612_/X sky130_fd_sc_hd__or4_1
X_4824_ _4831_/A _4824_/B _4824_/C vssd1 vssd1 vccd1 vccd1 _4961_/A sky130_fd_sc_hd__or3_2
XFILLER_21_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8592_ input3/X _8592_/D vssd1 vssd1 vccd1 vccd1 _8592_/Q sky130_fd_sc_hd__dfxtp_2
X_4755_ _4760_/A vssd1 vssd1 vccd1 vccd1 _5290_/A sky130_fd_sc_hd__clkbuf_4
X_7543_ _7543_/A _7543_/B vssd1 vssd1 vccd1 vccd1 _7543_/X sky130_fd_sc_hd__or2_1
X_7474_ _7474_/A _7474_/B vssd1 vssd1 vccd1 vccd1 _7474_/X sky130_fd_sc_hd__xor2_1
X_4686_ _4686_/A vssd1 vssd1 vccd1 vccd1 _5259_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6425_ _6425_/A vssd1 vssd1 vccd1 vccd1 _8670_/D sky130_fd_sc_hd__clkbuf_1
X_6356_ _6357_/A _6371_/B vssd1 vssd1 vccd1 vccd1 _6358_/A sky130_fd_sc_hd__and2_1
XFILLER_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5307_ _8635_/Q _8634_/Q _5306_/X _8636_/Q vssd1 vssd1 vccd1 vccd1 _5307_/X sky130_fd_sc_hd__a31o_1
X_8026_ _8116_/C _8115_/A vssd1 vssd1 vccd1 vccd1 _8026_/Y sky130_fd_sc_hd__nor2_1
X_6287_ _6287_/A _6287_/B vssd1 vssd1 vccd1 vccd1 _6290_/A sky130_fd_sc_hd__xnor2_1
XFILLER_102_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5238_ _5238_/A _5239_/B _5238_/C _5237_/Y vssd1 vssd1 vccd1 vccd1 _5238_/X sky130_fd_sc_hd__or4b_1
X_5169_ _5047_/D _5166_/X _5168_/X _5224_/C vssd1 vssd1 vccd1 vccd1 _5169_/X sky130_fd_sc_hd__o22a_1
XFILLER_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8928_ _8928_/A _4455_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[37] sky130_fd_sc_hd__ebufn_8
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8859_ _8859_/A _4374_/Y vssd1 vssd1 vccd1 vccd1 io_out[6] sky130_fd_sc_hd__ebufn_8
XFILLER_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4540_ _4831_/C _4849_/B _4822_/C vssd1 vssd1 vccd1 vccd1 _4861_/A sky130_fd_sc_hd__nand3b_4
XFILLER_7_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4471_ _4662_/A _4533_/B vssd1 vssd1 vccd1 vccd1 _4475_/C sky130_fd_sc_hd__nor2_1
X_7190_ _7190_/A _7190_/B vssd1 vssd1 vccd1 vccd1 _7208_/A sky130_fd_sc_hd__xnor2_1
XFILLER_99_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6210_ _6210_/A _6020_/A vssd1 vssd1 vccd1 vccd1 _6210_/X sky130_fd_sc_hd__or2b_1
X_6141_ _6303_/A _6141_/B vssd1 vssd1 vccd1 vccd1 _6300_/A sky130_fd_sc_hd__nand2_1
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6072_ _6072_/A _6072_/B vssd1 vssd1 vccd1 vccd1 _6103_/C sky130_fd_sc_hd__xor2_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5023_ _5023_/A vssd1 vssd1 vccd1 vccd1 _5190_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_65_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6974_ _6637_/A _6847_/A _6848_/A _6848_/B vssd1 vssd1 vccd1 vccd1 _7013_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_80_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8713_ input3/X _8713_/D vssd1 vssd1 vccd1 vccd1 _8713_/Q sky130_fd_sc_hd__dfxtp_1
X_5925_ _6277_/A _5951_/B vssd1 vssd1 vccd1 vccd1 _5926_/B sky130_fd_sc_hd__xor2_1
X_5856_ _5856_/A _5856_/B vssd1 vssd1 vccd1 vccd1 _5857_/B sky130_fd_sc_hd__or2_1
XFILLER_34_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8644_ input3/X _8644_/D vssd1 vssd1 vccd1 vccd1 _8644_/Q sky130_fd_sc_hd__dfxtp_1
X_4807_ _5180_/C _5253_/C vssd1 vssd1 vccd1 vccd1 _4899_/A sky130_fd_sc_hd__or2_1
X_8575_ input3/X _8575_/D vssd1 vssd1 vccd1 vccd1 _8575_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5787_ _5770_/A _5770_/B _5786_/X vssd1 vssd1 vccd1 vccd1 _5845_/A sky130_fd_sc_hd__a21oi_1
X_7526_ _7526_/A _7526_/B vssd1 vssd1 vccd1 vccd1 _7527_/B sky130_fd_sc_hd__nand2_1
X_4738_ _4802_/B vssd1 vssd1 vccd1 vccd1 _4850_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_7457_ _7458_/B _7458_/C _7458_/A vssd1 vssd1 vccd1 vccd1 _7459_/A sky130_fd_sc_hd__a21oi_1
X_4669_ _5045_/A vssd1 vssd1 vccd1 vccd1 _5235_/A sky130_fd_sc_hd__clkbuf_2
X_6408_ _8666_/Q _8665_/Q vssd1 vssd1 vccd1 vccd1 _6409_/C sky130_fd_sc_hd__nand2_1
X_7388_ _7388_/A _7388_/B _7388_/C vssd1 vssd1 vccd1 vccd1 _7409_/A sky130_fd_sc_hd__or3_1
X_6339_ _6329_/X _6338_/X _6334_/X _8656_/Q vssd1 vssd1 vccd1 vccd1 _8656_/D sky130_fd_sc_hd__o2bb2a_1
XFILLER_95_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8009_ _8019_/A _8009_/B _8009_/C vssd1 vssd1 vccd1 vccd1 _8019_/B sky130_fd_sc_hd__nand3_1
XFILLER_91_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5710_ _5768_/B _5710_/B vssd1 vssd1 vccd1 vccd1 _5861_/A sky130_fd_sc_hd__nand2_1
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6690_ _6718_/S _6724_/B _6689_/X vssd1 vssd1 vccd1 vccd1 _6691_/B sky130_fd_sc_hd__a21o_1
XFILLER_31_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5641_ _5641_/A vssd1 vssd1 vccd1 vccd1 _5642_/B sky130_fd_sc_hd__inv_2
X_8360_ _8360_/A _8360_/B vssd1 vssd1 vccd1 vccd1 _8365_/A sky130_fd_sc_hd__nand2_1
X_5572_ _6005_/A _6006_/A vssd1 vssd1 vccd1 vccd1 _5574_/B sky130_fd_sc_hd__nor2_1
X_8291_ _8368_/B _8291_/B vssd1 vssd1 vccd1 vccd1 _8295_/A sky130_fd_sc_hd__xor2_1
X_7311_ _7310_/A _7311_/B vssd1 vssd1 vccd1 vccd1 _7311_/X sky130_fd_sc_hd__and2b_1
X_4523_ _4727_/A vssd1 vssd1 vccd1 vccd1 _5149_/A sky130_fd_sc_hd__clkbuf_2
X_7242_ _7320_/A _7320_/B _7241_/Y vssd1 vssd1 vccd1 vccd1 _7268_/A sky130_fd_sc_hd__a21o_1
XFILLER_104_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4454_ _4456_/A vssd1 vssd1 vccd1 vccd1 _4454_/Y sky130_fd_sc_hd__inv_2
X_4385_ _4389_/A vssd1 vssd1 vccd1 vccd1 _4385_/Y sky130_fd_sc_hd__inv_2
X_7173_ _7173_/A _7188_/A vssd1 vssd1 vccd1 vccd1 _7272_/A sky130_fd_sc_hd__xor2_1
XFILLER_98_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6124_ _6125_/A _6125_/B vssd1 vssd1 vccd1 vccd1 _6124_/Y sky130_fd_sc_hd__nand2_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6055_ _6077_/A _6077_/B _6054_/Y vssd1 vssd1 vccd1 vccd1 _6057_/B sky130_fd_sc_hd__a21oi_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5006_ _5006_/A vssd1 vssd1 vccd1 vccd1 _5185_/C sky130_fd_sc_hd__clkbuf_2
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6957_ _6637_/A _6831_/B _7006_/A vssd1 vssd1 vccd1 vccd1 _7139_/A sky130_fd_sc_hd__mux2_1
X_8800__78 vssd1 vssd1 vccd1 vccd1 _8800__78/HI _8909_/A sky130_fd_sc_hd__conb_1
XFILLER_41_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6888_ _6868_/A _6868_/B _6870_/X vssd1 vssd1 vccd1 vccd1 _6888_/X sky130_fd_sc_hd__a21o_1
X_5908_ _5909_/A _6229_/A vssd1 vssd1 vccd1 vccd1 _6017_/B sky130_fd_sc_hd__nand2_1
X_8627_ input3/X _8627_/D vssd1 vssd1 vccd1 vccd1 _8627_/Q sky130_fd_sc_hd__dfxtp_1
X_5839_ _5920_/B _5920_/C vssd1 vssd1 vccd1 vccd1 _5840_/B sky130_fd_sc_hd__and2_1
X_8558_ _8566_/A _6427_/X _8557_/X vssd1 vssd1 vccd1 vccd1 _8723_/D sky130_fd_sc_hd__a21bo_1
XFILLER_14_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7509_ _7509_/A _7509_/B vssd1 vssd1 vccd1 vccd1 _7509_/Y sky130_fd_sc_hd__nor2_1
XFILLER_5_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8489_ _8490_/A _8490_/B _8490_/C vssd1 vssd1 vccd1 vccd1 _8489_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_89_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7860_ _7886_/A _7962_/B _7743_/B _7859_/Y vssd1 vssd1 vccd1 vccd1 _7867_/A sky130_fd_sc_hd__a31o_1
XFILLER_63_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6811_ _7160_/B _7031_/S vssd1 vssd1 vccd1 vccd1 _6812_/B sky130_fd_sc_hd__xor2_1
XFILLER_63_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7791_ _7800_/A _7904_/C vssd1 vssd1 vccd1 vccd1 _7792_/B sky130_fd_sc_hd__xnor2_1
XFILLER_50_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6742_ _7223_/B vssd1 vssd1 vccd1 vccd1 _7226_/B sky130_fd_sc_hd__clkbuf_2
X_6673_ _6673_/A vssd1 vssd1 vccd1 vccd1 _6769_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_8412_ _8412_/A _8412_/B vssd1 vssd1 vccd1 vccd1 _8412_/Y sky130_fd_sc_hd__nand2_1
X_5624_ _8650_/Q _6617_/A vssd1 vssd1 vccd1 vccd1 _5624_/X sky130_fd_sc_hd__and2b_1
X_8343_ _8343_/A _8343_/B vssd1 vssd1 vccd1 vccd1 _8377_/B sky130_fd_sc_hd__xnor2_1
X_5555_ _5554_/A _5554_/B _5553_/X vssd1 vssd1 vccd1 vccd1 _5556_/C sky130_fd_sc_hd__o21bai_1
X_8274_ _8201_/A _8201_/B _8202_/B _8202_/A vssd1 vssd1 vccd1 vccd1 _8297_/A sky130_fd_sc_hd__o2bb2a_1
X_4506_ _4831_/A vssd1 vssd1 vccd1 vccd1 _4849_/A sky130_fd_sc_hd__clkbuf_1
X_5486_ _5486_/A _5486_/B vssd1 vssd1 vccd1 vccd1 _5539_/A sky130_fd_sc_hd__xnor2_2
XFILLER_104_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7225_ _7230_/A _7434_/A vssd1 vssd1 vccd1 vccd1 _7307_/B sky130_fd_sc_hd__nor2_1
X_4437_ _4438_/A vssd1 vssd1 vccd1 vccd1 _4437_/Y sky130_fd_sc_hd__inv_2
X_7156_ _7156_/A _7156_/B vssd1 vssd1 vccd1 vccd1 _7157_/B sky130_fd_sc_hd__xnor2_2
X_4368_ _4370_/A vssd1 vssd1 vccd1 vccd1 _4368_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6107_ _6323_/C _6107_/B vssd1 vssd1 vccd1 vccd1 _6123_/B sky130_fd_sc_hd__or2_1
X_7087_ _7087_/A _7087_/B vssd1 vssd1 vccd1 vccd1 _7462_/B sky130_fd_sc_hd__xnor2_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6038_ _6038_/A _6038_/B _6038_/C vssd1 vssd1 vccd1 vccd1 _6060_/A sky130_fd_sc_hd__and3_1
XFILLER_46_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7989_ _8054_/A _8296_/A _8455_/A vssd1 vssd1 vccd1 vccd1 _8063_/A sky130_fd_sc_hd__a21bo_1
XFILLER_14_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8791__69 vssd1 vssd1 vccd1 vccd1 _8791__69/HI _8900_/A sky130_fd_sc_hd__conb_1
XFILLER_32_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5340_ _6475_/D _5342_/C _5374_/A vssd1 vssd1 vccd1 vccd1 _5340_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_5_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5271_ _5285_/A vssd1 vssd1 vccd1 vccd1 _5271_/X sky130_fd_sc_hd__clkbuf_2
X_7010_ _7010_/A _7010_/B _7010_/C vssd1 vssd1 vccd1 vccd1 _7011_/B sky130_fd_sc_hd__nand3_1
XFILLER_101_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7912_ _7912_/A _7912_/B vssd1 vssd1 vccd1 vccd1 _8455_/A sky130_fd_sc_hd__or2_4
XFILLER_24_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8892_ _8892_/A _4419_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[1] sky130_fd_sc_hd__ebufn_8
X_7843_ _7848_/A _8512_/A vssd1 vssd1 vccd1 vccd1 _7849_/A sky130_fd_sc_hd__nand2_1
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7774_ _7853_/B _8116_/B _7774_/C vssd1 vssd1 vccd1 vccd1 _7852_/B sky130_fd_sc_hd__and3_1
X_4986_ _5231_/D _4923_/X _5075_/B vssd1 vssd1 vccd1 vccd1 _4987_/D sky130_fd_sc_hd__o21a_1
X_6725_ _7293_/B _7246_/B _6676_/X _6692_/B _6724_/Y vssd1 vssd1 vccd1 vccd1 _6827_/A
+ sky130_fd_sc_hd__a32oi_4
XFILLER_51_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6656_ _6629_/A _6656_/B vssd1 vssd1 vccd1 vccd1 _6657_/A sky130_fd_sc_hd__and2b_1
XFILLER_31_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6587_ _7439_/A _6815_/B _6587_/C vssd1 vssd1 vccd1 vccd1 _6588_/C sky130_fd_sc_hd__and3_1
X_5607_ _5607_/A _5607_/B vssd1 vssd1 vccd1 vccd1 _5645_/B sky130_fd_sc_hd__nand2_1
X_8326_ _8326_/A _8326_/B vssd1 vssd1 vccd1 vccd1 _8334_/A sky130_fd_sc_hd__nor2_2
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5538_ _5558_/A _5516_/A _5551_/A vssd1 vssd1 vccd1 vccd1 _5540_/C sky130_fd_sc_hd__a21o_1
X_8257_ _8257_/A _8257_/B vssd1 vssd1 vccd1 vccd1 _8258_/B sky130_fd_sc_hd__xnor2_1
X_7208_ _7208_/A _7191_/A vssd1 vssd1 vccd1 vccd1 _7208_/X sky130_fd_sc_hd__or2b_1
X_5469_ _8660_/Q vssd1 vssd1 vccd1 vccd1 _6351_/A sky130_fd_sc_hd__inv_2
X_8188_ _8180_/A _8180_/B _8179_/A vssd1 vssd1 vccd1 vccd1 _8260_/A sky130_fd_sc_hd__o21ai_1
X_7139_ _7139_/A _7139_/B vssd1 vssd1 vccd1 vccd1 _7140_/B sky130_fd_sc_hd__xnor2_1
XFILLER_27_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4840_ _4865_/B _4960_/A vssd1 vssd1 vccd1 vccd1 _5101_/A sky130_fd_sc_hd__nor2_1
XFILLER_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4771_ _5263_/A _4775_/C vssd1 vssd1 vccd1 vccd1 _4772_/C sky130_fd_sc_hd__nand2_1
X_6510_ _6510_/A vssd1 vssd1 vccd1 vccd1 _8688_/D sky130_fd_sc_hd__clkbuf_1
X_7490_ _7490_/A _7490_/B vssd1 vssd1 vccd1 vccd1 _7490_/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6441_ _8676_/Q _6441_/B _6441_/C vssd1 vssd1 vccd1 vccd1 _6445_/B sky130_fd_sc_hd__and3_1
X_6372_ _6372_/A _6375_/B vssd1 vssd1 vccd1 vccd1 _6373_/B sky130_fd_sc_hd__nor2_1
X_8111_ _8205_/A _8111_/B _8111_/C vssd1 vssd1 vccd1 vccd1 _8126_/B sky130_fd_sc_hd__and3_1
X_5323_ _5323_/A vssd1 vssd1 vccd1 vccd1 _8626_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8042_ _8105_/B _8042_/B vssd1 vssd1 vccd1 vccd1 _8047_/A sky130_fd_sc_hd__xnor2_2
XFILLER_87_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5254_ _5143_/B _5118_/B _5252_/A _5248_/A _4885_/X vssd1 vssd1 vccd1 vccd1 _5256_/C
+ sky130_fd_sc_hd__a2111o_1
X_5185_ _5185_/A _5219_/B _5185_/C vssd1 vssd1 vccd1 vccd1 _5185_/X sky130_fd_sc_hd__or3_1
XFILLER_95_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8875_ _8875_/A _4393_/Y vssd1 vssd1 vccd1 vccd1 io_out[22] sky130_fd_sc_hd__ebufn_8
XFILLER_83_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7826_ _8207_/A _7839_/A _7777_/C _8116_/B vssd1 vssd1 vccd1 vccd1 _7841_/B sky130_fd_sc_hd__o211ai_2
XFILLER_51_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7757_ _7757_/A _7757_/B vssd1 vssd1 vccd1 vccd1 _7886_/C sky130_fd_sc_hd__xnor2_1
X_4969_ _5102_/C _4969_/B _4969_/C _5176_/C vssd1 vssd1 vccd1 vccd1 _4987_/C sky130_fd_sc_hd__or4_1
XFILLER_24_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6708_ _7223_/A _6806_/A vssd1 vssd1 vccd1 vccd1 _6765_/B sky130_fd_sc_hd__nor2_2
X_7688_ _8723_/Q _7688_/B vssd1 vssd1 vccd1 vccd1 _7747_/A sky130_fd_sc_hd__nor2_2
X_6639_ _6639_/A vssd1 vssd1 vccd1 vccd1 _6947_/A sky130_fd_sc_hd__buf_2
XFILLER_22_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8309_ _8302_/A _8384_/B _8437_/B _8287_/A vssd1 vssd1 vccd1 vccd1 _8310_/B sky130_fd_sc_hd__o22a_1
XFILLER_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8761__39 vssd1 vssd1 vccd1 vccd1 _8761__39/HI _8856_/A sky130_fd_sc_hd__conb_1
XFILLER_42_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6990_ _6853_/X _6894_/Y _6988_/X _6989_/Y vssd1 vssd1 vccd1 vccd1 _6995_/A sky130_fd_sc_hd__o211a_1
XFILLER_92_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5941_ _5941_/A _5941_/B vssd1 vssd1 vccd1 vccd1 _6074_/C sky130_fd_sc_hd__xor2_1
XFILLER_25_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5872_ _6205_/A _5873_/B vssd1 vssd1 vccd1 vccd1 _5991_/A sky130_fd_sc_hd__and2_1
X_8660_ input3/X _8660_/D vssd1 vssd1 vccd1 vccd1 _8660_/Q sky130_fd_sc_hd__dfxtp_1
X_7611_ _7611_/A _7611_/B _7611_/C vssd1 vssd1 vccd1 vccd1 _7622_/S sky130_fd_sc_hd__and3_1
X_4823_ _4823_/A _4823_/B vssd1 vssd1 vccd1 vccd1 _4898_/A sky130_fd_sc_hd__nor2_2
X_8591_ input3/X _8591_/D vssd1 vssd1 vccd1 vccd1 _8591_/Q sky130_fd_sc_hd__dfxtp_2
X_7542_ _7537_/A _7540_/A _7540_/Y _7541_/X vssd1 vssd1 vccd1 vccd1 _8704_/D sky130_fd_sc_hd__a211o_1
X_4754_ _4745_/A _4850_/B _5026_/A _4507_/X vssd1 vssd1 vccd1 vccd1 _4754_/X sky130_fd_sc_hd__a31o_1
X_7473_ _7449_/X _7473_/B vssd1 vssd1 vccd1 vccd1 _7474_/A sky130_fd_sc_hd__and2b_1
X_4685_ _5159_/A vssd1 vssd1 vccd1 vccd1 _4686_/A sky130_fd_sc_hd__clkbuf_2
X_6424_ _6430_/C _6424_/B _6461_/B vssd1 vssd1 vccd1 vccd1 _6425_/A sky130_fd_sc_hd__and3b_1
X_6355_ _5462_/B _5412_/X _5413_/X _6354_/Y vssd1 vssd1 vccd1 vccd1 _8660_/D sky130_fd_sc_hd__a22o_1
XFILLER_88_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5306_ _8631_/Q _8630_/Q _5304_/X _6475_/D _8633_/Q vssd1 vssd1 vccd1 vccd1 _5306_/X
+ sky130_fd_sc_hd__a311o_1
X_6286_ _6286_/A _6286_/B vssd1 vssd1 vccd1 vccd1 _6287_/B sky130_fd_sc_hd__xnor2_1
X_8025_ _8025_/A _8025_/B vssd1 vssd1 vccd1 vccd1 _8030_/A sky130_fd_sc_hd__nand2_1
X_5237_ _5227_/B _4823_/B _5072_/B vssd1 vssd1 vccd1 vccd1 _5237_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_75_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5168_ _5168_/A _5192_/B vssd1 vssd1 vccd1 vccd1 _5168_/X sky130_fd_sc_hd__or2_1
XFILLER_56_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5099_ _5139_/A _5097_/X _4937_/C _5098_/X _5040_/A vssd1 vssd1 vccd1 vccd1 _5099_/X
+ sky130_fd_sc_hd__o221a_1
X_8927_ _8927_/A _4454_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[36] sky130_fd_sc_hd__ebufn_8
XFILLER_83_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8858_ _8858_/A _4373_/Y vssd1 vssd1 vccd1 vccd1 io_out[5] sky130_fd_sc_hd__ebufn_8
XFILLER_24_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7809_ _7851_/A _7808_/C _7815_/A vssd1 vssd1 vccd1 vccd1 _7810_/B sky130_fd_sc_hd__o21ai_1
XFILLER_12_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8806__84 vssd1 vssd1 vccd1 vccd1 _8806__84/HI _8915_/A sky130_fd_sc_hd__conb_1
XFILLER_59_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4470_ _5226_/B _4705_/A vssd1 vssd1 vccd1 vccd1 _4533_/B sky130_fd_sc_hd__or2_1
X_6140_ _6140_/A _6140_/B _6140_/C vssd1 vssd1 vccd1 vccd1 _6141_/B sky130_fd_sc_hd__or3_1
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6071_ _6101_/A _6101_/B vssd1 vssd1 vccd1 vccd1 _6103_/B sky130_fd_sc_hd__and2_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5022_ _5003_/X _5192_/A _5014_/X _5021_/X vssd1 vssd1 vccd1 vccd1 _5022_/X sky130_fd_sc_hd__o31a_1
XFILLER_38_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6973_ _6973_/A _6885_/B vssd1 vssd1 vccd1 vccd1 _6982_/A sky130_fd_sc_hd__or2b_1
XFILLER_65_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8712_ input3/X _8712_/D vssd1 vssd1 vccd1 vccd1 _8712_/Q sky130_fd_sc_hd__dfxtp_1
X_5924_ _6185_/A _5828_/B _5869_/Y vssd1 vssd1 vccd1 vccd1 _5951_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5855_ _5856_/A _5856_/B vssd1 vssd1 vccd1 vccd1 _5857_/A sky130_fd_sc_hd__nand2_1
X_8643_ input3/X _8643_/D vssd1 vssd1 vccd1 vccd1 _8643_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4806_ _4861_/A _4897_/C vssd1 vssd1 vccd1 vccd1 _5253_/C sky130_fd_sc_hd__nor2_4
X_8574_ input3/X _8574_/D vssd1 vssd1 vccd1 vccd1 _8574_/Q sky130_fd_sc_hd__dfxtp_1
X_5786_ _5745_/A _5786_/B vssd1 vssd1 vccd1 vccd1 _5786_/X sky130_fd_sc_hd__and2b_1
X_7525_ _7525_/A _6711_/A vssd1 vssd1 vccd1 vccd1 _7526_/B sky130_fd_sc_hd__or2b_1
X_4737_ _4737_/A vssd1 vssd1 vccd1 vccd1 _8602_/D sky130_fd_sc_hd__clkbuf_1
X_7456_ _7456_/A _7456_/B vssd1 vssd1 vccd1 vccd1 _7458_/A sky130_fd_sc_hd__xnor2_1
X_4668_ _8592_/Q vssd1 vssd1 vccd1 vccd1 _5045_/A sky130_fd_sc_hd__inv_2
XFILLER_79_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6407_ _6461_/B vssd1 vssd1 vccd1 vccd1 _6409_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_103_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7387_ _7333_/Y _7382_/X _7381_/Y _7374_/X vssd1 vssd1 vccd1 vccd1 _7388_/C sky130_fd_sc_hd__o211a_1
X_4599_ _8575_/Q _4597_/A _4595_/X vssd1 vssd1 vccd1 vccd1 _4600_/B sky130_fd_sc_hd__o21ai_1
X_6338_ _6340_/S _6337_/X _6341_/A _6341_/B vssd1 vssd1 vccd1 vccd1 _6338_/X sky130_fd_sc_hd__a211o_1
XFILLER_103_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6269_ _6269_/A _6269_/B vssd1 vssd1 vccd1 vccd1 _6270_/B sky130_fd_sc_hd__or2_1
X_8008_ _8018_/A _8018_/B vssd1 vssd1 vccd1 vccd1 _8009_/C sky130_fd_sc_hd__xor2_1
XFILLER_57_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5640_ _5679_/A _5680_/A _5680_/B _5624_/X vssd1 vssd1 vccd1 vccd1 _5643_/A sky130_fd_sc_hd__a31o_2
XFILLER_31_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5571_ _5571_/A _5576_/B _5571_/C vssd1 vssd1 vccd1 vccd1 _5575_/A sky130_fd_sc_hd__nand3_1
X_8290_ _8290_/A _8290_/B vssd1 vssd1 vccd1 vccd1 _8291_/B sky130_fd_sc_hd__xnor2_1
X_7310_ _7310_/A _7311_/B vssd1 vssd1 vccd1 vccd1 _7332_/B sky130_fd_sc_hd__xnor2_1
X_4522_ _7708_/B vssd1 vssd1 vccd1 vccd1 _4727_/A sky130_fd_sc_hd__clkbuf_2
X_4453_ _4456_/A vssd1 vssd1 vccd1 vccd1 _4453_/Y sky130_fd_sc_hd__inv_2
X_7241_ _7241_/A _7241_/B vssd1 vssd1 vccd1 vccd1 _7241_/Y sky130_fd_sc_hd__nor2_1
XFILLER_7_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4384_ _4396_/A vssd1 vssd1 vccd1 vccd1 _4389_/A sky130_fd_sc_hd__clkbuf_4
X_7172_ _7172_/A _7172_/B vssd1 vssd1 vccd1 vccd1 _7188_/A sky130_fd_sc_hd__xor2_1
XFILLER_98_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6123_ _6123_/A _6123_/B vssd1 vssd1 vccd1 vccd1 _6142_/A sky130_fd_sc_hd__or2_2
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6054_ _6054_/A _6054_/B vssd1 vssd1 vccd1 vccd1 _6054_/Y sky130_fd_sc_hd__nor2_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5005_ _5005_/A vssd1 vssd1 vccd1 vccd1 _5182_/C sky130_fd_sc_hd__clkbuf_2
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8797__75 vssd1 vssd1 vccd1 vccd1 _8797__75/HI _8906_/A sky130_fd_sc_hd__conb_1
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6956_ _7417_/A _7219_/A _7226_/B vssd1 vssd1 vccd1 vccd1 _7010_/A sky130_fd_sc_hd__or3b_1
XFILLER_81_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5907_ _5907_/A _5907_/B vssd1 vssd1 vccd1 vccd1 _6229_/A sky130_fd_sc_hd__or2_2
X_6887_ _6887_/A _6887_/B vssd1 vssd1 vccd1 vccd1 _6968_/B sky130_fd_sc_hd__xor2_1
X_8626_ input3/X _8626_/D vssd1 vssd1 vccd1 vccd1 _8626_/Q sky130_fd_sc_hd__dfxtp_1
X_5838_ _5838_/A _5838_/B vssd1 vssd1 vccd1 vccd1 _5920_/C sky130_fd_sc_hd__or2_1
X_8557_ _8557_/A _8568_/A _8557_/C _8567_/S vssd1 vssd1 vccd1 vccd1 _8557_/X sky130_fd_sc_hd__or4_1
X_5769_ _5856_/A _5769_/B vssd1 vssd1 vccd1 vccd1 _5770_/B sky130_fd_sc_hd__nor2_1
X_7508_ _7508_/A _7508_/B vssd1 vssd1 vccd1 vccd1 _7509_/B sky130_fd_sc_hd__xnor2_1
X_8488_ _8488_/A _8488_/B vssd1 vssd1 vccd1 vccd1 _8490_/C sky130_fd_sc_hd__xor2_1
X_7439_ _7439_/A _7440_/B vssd1 vssd1 vccd1 vccd1 _7443_/B sky130_fd_sc_hd__xnor2_1
XFILLER_30_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6810_ _6947_/B vssd1 vssd1 vccd1 vccd1 _7031_/S sky130_fd_sc_hd__clkbuf_2
X_7790_ _7790_/A _8302_/A vssd1 vssd1 vccd1 vccd1 _7904_/C sky130_fd_sc_hd__nor2_1
X_6741_ _6806_/B vssd1 vssd1 vccd1 vccd1 _7223_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_50_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6672_ _7237_/B _7175_/B _7237_/C _7299_/A vssd1 vssd1 vccd1 vccd1 _6673_/A sky130_fd_sc_hd__or4b_1
X_8411_ _8412_/A _8412_/B _8409_/X vssd1 vssd1 vccd1 vccd1 _8471_/A sky130_fd_sc_hd__o21a_1
X_5623_ _5606_/A _5657_/B _5638_/B _5622_/X vssd1 vssd1 vccd1 vccd1 _5680_/B sky130_fd_sc_hd__a211o_1
X_8342_ _8342_/A _8342_/B vssd1 vssd1 vccd1 vccd1 _8343_/B sky130_fd_sc_hd__nor2_1
X_5554_ _5554_/A _5554_/B _5553_/X vssd1 vssd1 vccd1 vccd1 _5577_/B sky130_fd_sc_hd__or3b_1
X_8273_ _8258_/A _8258_/B _8272_/Y vssd1 vssd1 vccd1 vccd1 _8351_/B sky130_fd_sc_hd__a21o_1
X_4505_ _5607_/B vssd1 vssd1 vccd1 vccd1 _4831_/A sky130_fd_sc_hd__clkbuf_1
X_5485_ _5881_/A _5516_/A vssd1 vssd1 vccd1 vccd1 _5512_/A sky130_fd_sc_hd__nand2_1
X_7224_ _7226_/A _6869_/A _7195_/A _7222_/X _7229_/A vssd1 vssd1 vccd1 vccd1 _7434_/A
+ sky130_fd_sc_hd__o32a_2
X_4436_ _4438_/A vssd1 vssd1 vccd1 vccd1 _4436_/Y sky130_fd_sc_hd__inv_2
X_4367_ _4370_/A vssd1 vssd1 vccd1 vccd1 _4367_/Y sky130_fd_sc_hd__inv_2
XFILLER_104_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7155_ _7155_/A _7155_/B vssd1 vssd1 vccd1 vccd1 _7156_/B sky130_fd_sc_hd__xnor2_1
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6106_ _6106_/A _6106_/B vssd1 vssd1 vccd1 vccd1 _6310_/A sky130_fd_sc_hd__nor2_1
X_7086_ _7086_/A _7086_/B vssd1 vssd1 vccd1 vccd1 _7087_/B sky130_fd_sc_hd__xnor2_2
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6037_ _6082_/B _5574_/B _5575_/A _5574_/D vssd1 vssd1 vccd1 vccd1 _6038_/C sky130_fd_sc_hd__a22o_1
XFILLER_100_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7988_ _7988_/A _8152_/A vssd1 vssd1 vccd1 vccd1 _8054_/A sky130_fd_sc_hd__nand2_1
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6939_ _7044_/A _7044_/B _7044_/C _7044_/D vssd1 vssd1 vccd1 vccd1 _6939_/X sky130_fd_sc_hd__o22a_1
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8609_ input3/X _8609_/D vssd1 vssd1 vccd1 vccd1 _8609_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5270_ _5213_/X _5269_/Y _5290_/A vssd1 vssd1 vccd1 vccd1 _5285_/A sky130_fd_sc_hd__o21ai_4
XFILLER_99_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7911_ _7988_/A _7911_/B vssd1 vssd1 vccd1 vccd1 _7911_/Y sky130_fd_sc_hd__nand2_1
X_8767__45 vssd1 vssd1 vccd1 vccd1 _8767__45/HI _8862_/A sky130_fd_sc_hd__conb_1
XFILLER_83_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8891_ _8891_/A _4456_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[0] sky130_fd_sc_hd__ebufn_8
XFILLER_102_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7842_ _8508_/A _8508_/B _7842_/C vssd1 vssd1 vccd1 vccd1 _8512_/A sky130_fd_sc_hd__and3_1
XFILLER_24_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7773_ _7885_/A _8118_/A vssd1 vssd1 vccd1 vccd1 _7774_/C sky130_fd_sc_hd__nand2_1
X_4985_ _5172_/A _4985_/B vssd1 vssd1 vccd1 vccd1 _5167_/B sky130_fd_sc_hd__or2_1
XFILLER_23_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6724_ _6724_/A _6724_/B vssd1 vssd1 vccd1 vccd1 _6724_/Y sky130_fd_sc_hd__nand2_1
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6655_ _6697_/A vssd1 vssd1 vccd1 vccd1 _7249_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6586_ _6580_/B _7236_/A _7297_/A vssd1 vssd1 vccd1 vccd1 _6587_/C sky130_fd_sc_hd__o21ai_1
X_5606_ _5606_/A vssd1 vssd1 vccd1 vccd1 _5657_/A sky130_fd_sc_hd__clkbuf_2
X_8325_ _8229_/A _8334_/B _7964_/X vssd1 vssd1 vccd1 vccd1 _8392_/A sky130_fd_sc_hd__a21o_1
X_5537_ _5724_/B _5724_/C vssd1 vssd1 vccd1 vccd1 _5540_/B sky130_fd_sc_hd__and2_1
X_8256_ _8256_/A _8256_/B vssd1 vssd1 vccd1 vccd1 _8257_/B sky130_fd_sc_hd__nand2_1
XFILLER_11_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7207_ _7259_/A _7207_/B vssd1 vssd1 vccd1 vccd1 _7278_/B sky130_fd_sc_hd__xnor2_1
XFILLER_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5468_ _5468_/A _5468_/B vssd1 vssd1 vccd1 vccd1 _5477_/B sky130_fd_sc_hd__nor2_2
X_8187_ _8185_/Y _8183_/B _8186_/X vssd1 vssd1 vccd1 vccd1 _8428_/A sky130_fd_sc_hd__a21boi_1
X_5399_ _8646_/Q vssd1 vssd1 vccd1 vccd1 _5421_/B sky130_fd_sc_hd__inv_2
X_4419_ _4420_/A vssd1 vssd1 vccd1 vccd1 _4419_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7138_ _7220_/A _7137_/B _7137_/X _6876_/A _6806_/A vssd1 vssd1 vccd1 vccd1 _7139_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_86_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7069_ _7101_/D _7069_/B _7069_/C vssd1 vssd1 vccd1 vccd1 _7072_/A sky130_fd_sc_hd__nand3_1
XFILLER_100_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4770_ _5263_/A _4775_/C vssd1 vssd1 vccd1 vccd1 _4772_/B sky130_fd_sc_hd__or2_1
X_6440_ _6441_/B _6441_/C _6439_/Y vssd1 vssd1 vccd1 vccd1 _8675_/D sky130_fd_sc_hd__a21oi_1
X_6371_ _6371_/A _6371_/B vssd1 vssd1 vccd1 vccd1 _6375_/B sky130_fd_sc_hd__nor2_1
X_8110_ _8321_/A _8031_/B _8109_/X vssd1 vssd1 vccd1 vccd1 _8214_/A sky130_fd_sc_hd__a21bo_1
X_5322_ _5324_/B _5354_/B _5322_/C vssd1 vssd1 vccd1 vccd1 _5323_/A sky130_fd_sc_hd__and3b_1
X_8041_ _8041_/A _8041_/B vssd1 vssd1 vccd1 vccd1 _8042_/B sky130_fd_sc_hd__xnor2_1
X_5253_ _5253_/A _5253_/B _5253_/C _5237_/Y vssd1 vssd1 vccd1 vccd1 _5253_/X sky130_fd_sc_hd__or4b_1
XFILLER_87_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5184_ _5219_/A _5214_/C _5181_/X _5182_/X _5183_/X vssd1 vssd1 vccd1 vccd1 _5184_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_56_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8874_ _8874_/A _4392_/Y vssd1 vssd1 vccd1 vccd1 io_out[21] sky130_fd_sc_hd__ebufn_8
XFILLER_71_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7825_ _8317_/A _7886_/A vssd1 vssd1 vccd1 vccd1 _7839_/A sky130_fd_sc_hd__nor2_1
XFILLER_51_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7756_ _7823_/A _8111_/B _8111_/C vssd1 vssd1 vccd1 vccd1 _7757_/B sky130_fd_sc_hd__and3_1
XFILLER_11_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4968_ _5231_/D _5009_/B _4923_/X _4657_/A vssd1 vssd1 vccd1 vccd1 _4970_/C sky130_fd_sc_hd__o31a_1
X_6707_ _6844_/A vssd1 vssd1 vccd1 vccd1 _7223_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7687_ _7687_/A _7687_/B vssd1 vssd1 vccd1 vccd1 _7814_/A sky130_fd_sc_hd__xnor2_1
X_4899_ _4899_/A _5153_/B vssd1 vssd1 vccd1 vccd1 _5074_/B sky130_fd_sc_hd__or2_2
X_6638_ _7175_/A vssd1 vssd1 vccd1 vccd1 _7418_/A sky130_fd_sc_hd__clkbuf_2
X_8308_ _8308_/A _8363_/B vssd1 vssd1 vccd1 vccd1 _8437_/B sky130_fd_sc_hd__xor2_1
X_6569_ _7245_/A vssd1 vssd1 vccd1 vccd1 _7297_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_3_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8239_ _8239_/A _8239_/B vssd1 vssd1 vccd1 vccd1 _8299_/B sky130_fd_sc_hd__xor2_2
XFILLER_59_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5940_ _5943_/A _5943_/B vssd1 vssd1 vccd1 vccd1 _5941_/B sky130_fd_sc_hd__xor2_1
XFILLER_92_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8737__15 vssd1 vssd1 vccd1 vccd1 _8737__15/HI _8832_/A sky130_fd_sc_hd__conb_1
XFILLER_33_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7610_ _7611_/A _7611_/B _7611_/C vssd1 vssd1 vccd1 vccd1 _7612_/C sky130_fd_sc_hd__a21oi_1
X_5871_ _6203_/A _5869_/Y _5870_/Y vssd1 vssd1 vccd1 vccd1 _5873_/B sky130_fd_sc_hd__a21oi_1
XFILLER_61_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4822_ _4822_/A _4849_/B _4822_/C vssd1 vssd1 vccd1 vccd1 _4823_/B sky130_fd_sc_hd__and3_2
X_8590_ input3/X _8590_/D vssd1 vssd1 vccd1 vccd1 _8590_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7541_ _8557_/A vssd1 vssd1 vccd1 vccd1 _7541_/X sky130_fd_sc_hd__buf_2
X_4753_ _4842_/C vssd1 vssd1 vccd1 vccd1 _5026_/A sky130_fd_sc_hd__clkbuf_2
X_7472_ _7494_/A _7496_/A vssd1 vssd1 vccd1 vccd1 _7505_/B sky130_fd_sc_hd__xnor2_1
X_4684_ _4684_/A vssd1 vssd1 vccd1 vccd1 _8593_/D sky130_fd_sc_hd__clkbuf_1
X_6423_ _8668_/Q _6397_/D _6416_/B _8670_/Q vssd1 vssd1 vccd1 vccd1 _6424_/B sky130_fd_sc_hd__a31o_1
X_6354_ _6354_/A _6354_/B vssd1 vssd1 vccd1 vccd1 _6354_/Y sky130_fd_sc_hd__xnor2_1
X_5305_ _8632_/Q vssd1 vssd1 vccd1 vccd1 _6475_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6285_ _6285_/A _6285_/B vssd1 vssd1 vccd1 vccd1 _6286_/B sky130_fd_sc_hd__xor2_1
XFILLER_88_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8024_ _8134_/B vssd1 vssd1 vccd1 vccd1 _8031_/A sky130_fd_sc_hd__buf_2
X_5236_ _5029_/B _5151_/A _5235_/X _5245_/B _5143_/B vssd1 vssd1 vccd1 vccd1 _5238_/C
+ sky130_fd_sc_hd__o32a_1
XFILLER_84_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5167_ _5243_/C _5167_/B _5193_/D vssd1 vssd1 vccd1 vccd1 _5192_/B sky130_fd_sc_hd__or3_1
XFILLER_83_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5098_ _5214_/A _5098_/B _5243_/C _5098_/D vssd1 vssd1 vccd1 vccd1 _5098_/X sky130_fd_sc_hd__or4_1
XFILLER_29_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8926_ _8926_/A _4453_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[35] sky130_fd_sc_hd__ebufn_8
XFILLER_83_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8857_ _8857_/A _4370_/Y vssd1 vssd1 vccd1 vccd1 io_out[4] sky130_fd_sc_hd__ebufn_8
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7808_ _7815_/A _7851_/A _7808_/C vssd1 vssd1 vccd1 vccd1 _7942_/A sky130_fd_sc_hd__or3_1
XFILLER_52_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7739_ _7739_/A _7764_/A vssd1 vssd1 vccd1 vccd1 _7758_/A sky130_fd_sc_hd__nand2_1
XFILLER_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6070_ _6070_/A _6070_/B vssd1 vssd1 vccd1 vccd1 _6101_/B sky130_fd_sc_hd__xnor2_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5021_ _5105_/A _5168_/A _5018_/X _5020_/X vssd1 vssd1 vccd1 vccd1 _5021_/X sky130_fd_sc_hd__a211o_1
XFILLER_38_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6972_ _7202_/A vssd1 vssd1 vccd1 vccd1 _7205_/A sky130_fd_sc_hd__clkinv_2
XFILLER_93_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8711_ input3/X _8711_/D vssd1 vssd1 vccd1 vccd1 _8711_/Q sky130_fd_sc_hd__dfxtp_1
X_5923_ _6323_/D _5923_/B vssd1 vssd1 vccd1 vccd1 _6270_/A sky130_fd_sc_hd__nand2_1
X_5854_ _5937_/B _5854_/B vssd1 vssd1 vccd1 vccd1 _5856_/B sky130_fd_sc_hd__xnor2_1
X_8642_ input3/X _8642_/D vssd1 vssd1 vccd1 vccd1 _8642_/Q sky130_fd_sc_hd__dfxtp_1
X_4805_ _4860_/A _4908_/A vssd1 vssd1 vccd1 vccd1 _5180_/C sky130_fd_sc_hd__nor2_2
X_8573_ input3/X _8573_/D vssd1 vssd1 vccd1 vccd1 _8573_/Q sky130_fd_sc_hd__dfxtp_1
X_7524_ _7522_/A _7522_/B _7520_/A vssd1 vssd1 vccd1 vccd1 _7527_/A sky130_fd_sc_hd__a21oi_1
X_5785_ _6032_/A _6032_/B _5784_/X vssd1 vssd1 vccd1 vccd1 _5862_/A sky130_fd_sc_hd__a21o_1
X_4736_ _4733_/Y _7503_/A _4736_/C vssd1 vssd1 vccd1 vccd1 _4737_/A sky130_fd_sc_hd__and3b_1
X_7455_ _7456_/A _7455_/B vssd1 vssd1 vccd1 vccd1 _7458_/C sky130_fd_sc_hd__nand2_1
X_4667_ _5176_/A vssd1 vssd1 vccd1 vccd1 _5243_/A sky130_fd_sc_hd__clkbuf_2
X_7386_ _7380_/A _7384_/Y _7385_/Y vssd1 vssd1 vccd1 vccd1 _7388_/B sky130_fd_sc_hd__o21a_1
X_6406_ _6406_/A _6406_/B vssd1 vssd1 vccd1 vccd1 _6461_/B sky130_fd_sc_hd__and2_1
XFILLER_1_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4598_ _8574_/Q _8575_/Q _4598_/C vssd1 vssd1 vccd1 vccd1 _4604_/C sky130_fd_sc_hd__and3_1
X_6337_ _6337_/A _6336_/A vssd1 vssd1 vccd1 vccd1 _6337_/X sky130_fd_sc_hd__or2b_1
XFILLER_88_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6268_ _6232_/A _6233_/A _6232_/B vssd1 vssd1 vccd1 vccd1 _6271_/A sky130_fd_sc_hd__o21ba_1
X_8007_ _8083_/A _8006_/Y _7985_/C _7922_/B vssd1 vssd1 vccd1 vccd1 _8018_/B sky130_fd_sc_hd__a2bb2o_1
X_5219_ _5219_/A _5219_/B _5219_/C _5219_/D vssd1 vssd1 vccd1 vccd1 _5219_/X sky130_fd_sc_hd__or4_1
X_6199_ _6199_/A _6199_/B vssd1 vssd1 vccd1 vccd1 _6199_/Y sky130_fd_sc_hd__nand2_1
XFILLER_28_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8909_ _8909_/A _4432_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[18] sky130_fd_sc_hd__ebufn_8
XFILLER_12_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5570_ _5569_/A _5569_/B _5568_/X vssd1 vssd1 vccd1 vccd1 _5571_/C sky130_fd_sc_hd__o21bai_1
X_4521_ _8595_/Q vssd1 vssd1 vccd1 vccd1 _7708_/B sky130_fd_sc_hd__buf_2
X_4452_ _4456_/A vssd1 vssd1 vccd1 vccd1 _4452_/Y sky130_fd_sc_hd__inv_2
X_7240_ _7241_/A _7241_/B vssd1 vssd1 vccd1 vccd1 _7320_/B sky130_fd_sc_hd__xor2_1
XFILLER_104_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7171_ _7262_/A _7262_/B _7262_/C _7162_/B _7266_/A vssd1 vssd1 vccd1 vccd1 _7173_/A
+ sky130_fd_sc_hd__a32o_1
X_4383_ _4383_/A vssd1 vssd1 vccd1 vccd1 _4383_/Y sky130_fd_sc_hd__inv_2
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6122_ _6135_/B _6122_/B vssd1 vssd1 vccd1 vccd1 _6131_/A sky130_fd_sc_hd__nand2_1
X_6053_ _6053_/A _6053_/B vssd1 vssd1 vccd1 vccd1 _6077_/B sky130_fd_sc_hd__xnor2_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5004_ _5245_/C _5240_/C _5004_/C vssd1 vssd1 vccd1 vccd1 _5192_/A sky130_fd_sc_hd__or3_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6955_ _7223_/A vssd1 vssd1 vccd1 vccd1 _7417_/A sky130_fd_sc_hd__clkbuf_2
X_5906_ _5906_/A _6014_/B vssd1 vssd1 vccd1 vccd1 _5909_/A sky130_fd_sc_hd__xnor2_1
X_6886_ _6886_/A _6886_/B vssd1 vssd1 vccd1 vccd1 _6887_/B sky130_fd_sc_hd__xnor2_1
XFILLER_34_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8625_ input3/X _8625_/D vssd1 vssd1 vccd1 vccd1 _8625_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5837_ _5838_/A _6205_/A vssd1 vssd1 vccd1 vccd1 _5920_/B sky130_fd_sc_hd__nand2_1
XFILLER_22_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8556_ _8556_/A _8556_/B _8556_/C vssd1 vssd1 vccd1 vccd1 _8567_/S sky130_fd_sc_hd__and3_1
X_5768_ _5768_/A _5768_/B _5768_/C vssd1 vssd1 vccd1 vccd1 _5769_/B sky130_fd_sc_hd__and3_1
X_8487_ _8487_/A _8487_/B vssd1 vssd1 vccd1 vccd1 _8488_/B sky130_fd_sc_hd__xnor2_1
X_7507_ _7503_/X _8697_/Q _7498_/Y _7506_/X vssd1 vssd1 vccd1 vccd1 _8697_/D sky130_fd_sc_hd__o22a_1
XFILLER_5_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4719_ _7753_/A vssd1 vssd1 vccd1 vccd1 _5265_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7438_ _7438_/A _7438_/B vssd1 vssd1 vccd1 vccd1 _7440_/B sky130_fd_sc_hd__xor2_1
X_5699_ _5699_/A _5699_/B vssd1 vssd1 vccd1 vccd1 _6040_/A sky130_fd_sc_hd__xnor2_1
XFILLER_30_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7369_ _7296_/B _7296_/C _7296_/A vssd1 vssd1 vccd1 vccd1 _7398_/B sky130_fd_sc_hd__o21ai_1
XFILLER_103_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6740_ _7030_/B _7301_/A vssd1 vssd1 vccd1 vccd1 _6868_/A sky130_fd_sc_hd__nand2_1
X_6671_ _6671_/A _6671_/B vssd1 vssd1 vccd1 vccd1 _7299_/A sky130_fd_sc_hd__nor2_1
XFILLER_31_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8410_ _8410_/A _8410_/B _8410_/C vssd1 vssd1 vccd1 vccd1 _8412_/B sky130_fd_sc_hd__and3_1
X_5622_ _8648_/Q _7631_/B vssd1 vssd1 vccd1 vccd1 _5622_/X sky130_fd_sc_hd__and2b_1
X_8341_ _8341_/A _8341_/B _8341_/C vssd1 vssd1 vccd1 vccd1 _8342_/B sky130_fd_sc_hd__and3_1
X_5553_ _5553_/A _5553_/B vssd1 vssd1 vccd1 vccd1 _5553_/X sky130_fd_sc_hd__xor2_1
X_4504_ _7627_/B vssd1 vssd1 vccd1 vccd1 _5607_/B sky130_fd_sc_hd__clkbuf_2
X_8272_ _8272_/A _8272_/B vssd1 vssd1 vccd1 vccd1 _8272_/Y sky130_fd_sc_hd__nor2_1
X_5484_ _5520_/A _5520_/B vssd1 vssd1 vccd1 vccd1 _5516_/A sky130_fd_sc_hd__xor2_1
X_7223_ _7223_/A _7223_/B vssd1 vssd1 vccd1 vccd1 _7229_/A sky130_fd_sc_hd__or2_1
X_4435_ _4438_/A vssd1 vssd1 vccd1 vccd1 _4435_/Y sky130_fd_sc_hd__inv_2
X_4366_ _4370_/A vssd1 vssd1 vccd1 vccd1 _4366_/Y sky130_fd_sc_hd__inv_2
X_7154_ _7084_/A _7083_/B _7083_/A vssd1 vssd1 vccd1 vccd1 _7155_/B sky130_fd_sc_hd__o21bai_1
XFILLER_98_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6105_ _6167_/A _6104_/B _6102_/X vssd1 vssd1 vccd1 vccd1 _6106_/B sky130_fd_sc_hd__a21boi_1
X_7085_ _7147_/A _7147_/B vssd1 vssd1 vccd1 vccd1 _7086_/B sky130_fd_sc_hd__xnor2_2
XFILLER_58_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6036_ _6081_/A _6081_/B vssd1 vssd1 vccd1 vccd1 _6038_/B sky130_fd_sc_hd__nor2_1
XFILLER_27_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7987_ _7784_/B _7786_/B _7908_/X vssd1 vssd1 vccd1 vccd1 _8152_/A sky130_fd_sc_hd__a21oi_4
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6938_ _7044_/A _7044_/B _7044_/C _7044_/D vssd1 vssd1 vccd1 vccd1 _6938_/Y sky130_fd_sc_hd__nor4_2
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6869_ _6869_/A vssd1 vssd1 vccd1 vccd1 _7137_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_8608_ input3/X _8608_/D vssd1 vssd1 vccd1 vccd1 _8608_/Q sky130_fd_sc_hd__dfxtp_2
X_8539_ _8539_/A _8539_/B vssd1 vssd1 vccd1 vccd1 _8540_/B sky130_fd_sc_hd__nor2_1
XFILLER_10_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8890_ _8890_/A _4422_/Y vssd1 vssd1 vccd1 vccd1 io_out[37] sky130_fd_sc_hd__ebufn_8
XFILLER_83_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7910_ _7912_/B vssd1 vssd1 vccd1 vccd1 _8296_/A sky130_fd_sc_hd__buf_2
X_7841_ _7841_/A _7841_/B vssd1 vssd1 vccd1 vccd1 _7842_/C sky130_fd_sc_hd__xor2_1
XFILLER_48_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7772_ _7772_/A _7772_/B vssd1 vssd1 vccd1 vccd1 _7775_/A sky130_fd_sc_hd__xnor2_1
XFILLER_51_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4984_ _5135_/A vssd1 vssd1 vccd1 vccd1 _5219_/A sky130_fd_sc_hd__buf_2
X_6723_ _6723_/A vssd1 vssd1 vccd1 vccd1 _7246_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_23_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6654_ _7176_/B _7176_/C vssd1 vssd1 vccd1 vccd1 _6697_/A sky130_fd_sc_hd__and2_1
X_5605_ _7627_/B _8647_/Q vssd1 vssd1 vccd1 vccd1 _5606_/A sky130_fd_sc_hd__or2b_1
X_6585_ _7193_/A vssd1 vssd1 vccd1 vccd1 _7236_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_11_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8324_ _8324_/A _8324_/B vssd1 vssd1 vccd1 vccd1 _8341_/A sky130_fd_sc_hd__or2_1
X_5536_ _5558_/A _5551_/A _5492_/B _5560_/A vssd1 vssd1 vccd1 vccd1 _5542_/A sky130_fd_sc_hd__a22o_1
X_8255_ _8255_/A _8255_/B vssd1 vssd1 vccd1 vccd1 _8257_/A sky130_fd_sc_hd__nor2_1
X_5467_ _7699_/B _8661_/Q vssd1 vssd1 vccd1 vccd1 _5468_/B sky130_fd_sc_hd__and2b_1
X_7206_ _7206_/A _7206_/B vssd1 vssd1 vccd1 vccd1 _7207_/B sky130_fd_sc_hd__xor2_2
X_4418_ _4420_/A vssd1 vssd1 vccd1 vccd1 _4418_/Y sky130_fd_sc_hd__inv_2
X_8186_ _8186_/A _8182_/B vssd1 vssd1 vccd1 vccd1 _8186_/X sky130_fd_sc_hd__or2b_1
X_5398_ _5441_/A _5447_/A _5397_/X _8653_/Q vssd1 vssd1 vccd1 vccd1 _5398_/Y sky130_fd_sc_hd__a31oi_1
X_4349_ _4352_/A vssd1 vssd1 vccd1 vccd1 _4349_/Y sky130_fd_sc_hd__inv_2
X_7137_ _7226_/A _7137_/B vssd1 vssd1 vccd1 vccd1 _7137_/X sky130_fd_sc_hd__or2_1
XFILLER_100_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7068_ _7068_/A _7068_/B vssd1 vssd1 vccd1 vccd1 _7069_/C sky130_fd_sc_hd__xor2_1
XFILLER_74_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6019_ _6019_/A _6019_/B vssd1 vssd1 vccd1 vccd1 _6210_/A sky130_fd_sc_hd__xnor2_1
XFILLER_39_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6370_ _6371_/A _6371_/B vssd1 vssd1 vccd1 vccd1 _6372_/A sky130_fd_sc_hd__and2_1
X_5321_ _8625_/Q _8624_/Q _8626_/Q vssd1 vssd1 vccd1 vccd1 _5322_/C sky130_fd_sc_hd__a21o_1
X_8040_ _8040_/A _8040_/B vssd1 vssd1 vccd1 vccd1 _8041_/B sky130_fd_sc_hd__xnor2_1
XFILLER_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5252_ _5252_/A _5252_/B vssd1 vssd1 vccd1 vccd1 _5252_/X sky130_fd_sc_hd__or2_1
X_5183_ _5173_/D _5176_/D _5183_/S vssd1 vssd1 vccd1 vccd1 _5183_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8873_ _8873_/A _4391_/Y vssd1 vssd1 vccd1 vccd1 io_out[20] sky130_fd_sc_hd__ebufn_8
XFILLER_36_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7824_ _7884_/A vssd1 vssd1 vccd1 vccd1 _8317_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_36_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7755_ _7766_/A _7766_/C _7766_/B vssd1 vssd1 vccd1 vccd1 _8111_/C sky130_fd_sc_hd__a21o_1
XFILLER_51_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4967_ _5086_/A _5165_/C vssd1 vssd1 vccd1 vccd1 _5231_/D sky130_fd_sc_hd__or2_2
X_6706_ _7172_/A _7172_/B vssd1 vssd1 vccd1 vccd1 _6734_/B sky130_fd_sc_hd__or2b_1
X_7686_ _7687_/A _7687_/B _7685_/X _7664_/X vssd1 vssd1 vccd1 vccd1 _7812_/A sky130_fd_sc_hd__o2bb2a_1
X_4898_ _4898_/A _4898_/B vssd1 vssd1 vccd1 vccd1 _5153_/B sky130_fd_sc_hd__nor2_4
X_6637_ _6637_/A _6772_/A vssd1 vssd1 vccd1 vccd1 _6831_/B sky130_fd_sc_hd__nand2_2
X_6568_ _6591_/A _6591_/B vssd1 vssd1 vccd1 vccd1 _7245_/A sky130_fd_sc_hd__and2_1
X_8307_ _8384_/B _8385_/B vssd1 vssd1 vccd1 vccd1 _8363_/B sky130_fd_sc_hd__and2_1
X_5519_ _5896_/A _5794_/B _5794_/C vssd1 vssd1 vccd1 vccd1 _5906_/A sky130_fd_sc_hd__nand3_4
X_6499_ _6526_/B vssd1 vssd1 vccd1 vccd1 _6531_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_8238_ _8238_/A _8238_/B vssd1 vssd1 vccd1 vccd1 _8239_/B sky130_fd_sc_hd__xnor2_2
X_8169_ _8293_/A _8169_/B vssd1 vssd1 vccd1 vccd1 _8172_/B sky130_fd_sc_hd__and2_1
XFILLER_78_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5870_ _5983_/B _5870_/B vssd1 vssd1 vccd1 vccd1 _5870_/Y sky130_fd_sc_hd__nor2_1
XFILLER_18_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4821_ _4930_/A vssd1 vssd1 vccd1 vccd1 _4823_/A sky130_fd_sc_hd__inv_2
XFILLER_61_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7540_ _7540_/A _7540_/B vssd1 vssd1 vccd1 vccd1 _7540_/Y sky130_fd_sc_hd__nor2_1
X_4752_ _4752_/A vssd1 vssd1 vccd1 vccd1 _4856_/A sky130_fd_sc_hd__buf_2
XFILLER_21_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7471_ _7495_/A _7495_/B vssd1 vssd1 vccd1 vccd1 _7496_/A sky130_fd_sc_hd__nor2_1
X_4683_ _4717_/A _4683_/B _4707_/A vssd1 vssd1 vccd1 vccd1 _4684_/A sky130_fd_sc_hd__and3_1
X_6422_ _8669_/Q _8670_/Q _6422_/C vssd1 vssd1 vccd1 vccd1 _6430_/C sky130_fd_sc_hd__and3_1
X_6353_ _6343_/S _6348_/B _6347_/A vssd1 vssd1 vccd1 vccd1 _6354_/B sky130_fd_sc_hd__o21a_1
X_5304_ _8627_/Q _8626_/Q _6478_/A _6475_/B _8629_/Q vssd1 vssd1 vccd1 vccd1 _5304_/X
+ sky130_fd_sc_hd__a311o_1
X_6284_ _6203_/A _5986_/A _6284_/S vssd1 vssd1 vccd1 vccd1 _6285_/B sky130_fd_sc_hd__mux2_1
XFILLER_88_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8023_ _8023_/A _8023_/B vssd1 vssd1 vccd1 vccd1 _8107_/A sky130_fd_sc_hd__nand2_1
X_5235_ _5235_/A _5243_/B _5252_/A vssd1 vssd1 vccd1 vccd1 _5235_/X sky130_fd_sc_hd__or3_1
XFILLER_96_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5166_ _5166_/A _5166_/B _5231_/D _5166_/D vssd1 vssd1 vccd1 vccd1 _5166_/X sky130_fd_sc_hd__or4_1
XFILLER_68_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5097_ _4731_/A _5091_/X _5096_/X vssd1 vssd1 vccd1 vccd1 _5097_/X sky130_fd_sc_hd__o21a_1
X_8925_ _8925_/A _4452_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[34] sky130_fd_sc_hd__ebufn_8
XFILLER_17_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8856_ _8856_/A _4369_/Y vssd1 vssd1 vccd1 vccd1 io_out[3] sky130_fd_sc_hd__ebufn_8
X_7807_ _7807_/A _7807_/B vssd1 vssd1 vccd1 vccd1 _7808_/C sky130_fd_sc_hd__and2_1
XFILLER_52_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5999_ _6000_/A _6000_/B vssd1 vssd1 vccd1 vccd1 _6001_/A sky130_fd_sc_hd__or2_1
X_7738_ _7864_/B vssd1 vssd1 vccd1 vccd1 _7764_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7669_ _7819_/A _7819_/B vssd1 vssd1 vccd1 vccd1 _7820_/A sky130_fd_sc_hd__nor2_1
XFILLER_79_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5020_ _5135_/A _5239_/B _5215_/C _5047_/B vssd1 vssd1 vccd1 vccd1 _5020_/X sky130_fd_sc_hd__or4_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6971_ _6851_/A _6851_/B _6970_/X vssd1 vssd1 vccd1 vccd1 _6996_/B sky130_fd_sc_hd__a21o_1
XFILLER_80_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8710_ input3/X _8710_/D vssd1 vssd1 vccd1 vccd1 _8710_/Q sky130_fd_sc_hd__dfxtp_1
X_5922_ _5922_/A vssd1 vssd1 vccd1 vccd1 _6323_/D sky130_fd_sc_hd__buf_2
XFILLER_46_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5853_ _5777_/A _5777_/C _5777_/B vssd1 vssd1 vccd1 vccd1 _5854_/B sky130_fd_sc_hd__a21boi_1
X_8641_ input3/X _8641_/D vssd1 vssd1 vccd1 vccd1 _8641_/Q sky130_fd_sc_hd__dfxtp_1
X_4804_ _4829_/A vssd1 vssd1 vccd1 vccd1 _4908_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_21_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8572_ input3/X _8572_/D vssd1 vssd1 vccd1 vccd1 _8572_/Q sky130_fd_sc_hd__dfxtp_1
X_5784_ _5771_/A _5784_/B vssd1 vssd1 vccd1 vccd1 _5784_/X sky130_fd_sc_hd__and2b_1
X_7523_ _7518_/B _6511_/X _6513_/A _7522_/X vssd1 vssd1 vccd1 vccd1 _8701_/D sky130_fd_sc_hd__a22o_1
XFILLER_9_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4735_ _4909_/A _4739_/B vssd1 vssd1 vccd1 vccd1 _4736_/C sky130_fd_sc_hd__nand2_1
XFILLER_21_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7454_ _7454_/A _7363_/B vssd1 vssd1 vccd1 vccd1 _7458_/B sky130_fd_sc_hd__or2b_1
X_4666_ _5068_/A vssd1 vssd1 vccd1 vccd1 _5176_/A sky130_fd_sc_hd__clkbuf_2
X_7385_ _7385_/A _7385_/B vssd1 vssd1 vccd1 vccd1 _7385_/Y sky130_fd_sc_hd__nand2_1
X_4597_ _4597_/A _4597_/B vssd1 vssd1 vccd1 vccd1 _8574_/D sky130_fd_sc_hd__nor2_1
X_6405_ _6405_/A vssd1 vssd1 vccd1 vccd1 _8665_/D sky130_fd_sc_hd__clkbuf_1
X_6336_ _6336_/A _6337_/A vssd1 vssd1 vccd1 vccd1 _6340_/S sky130_fd_sc_hd__or2b_1
XFILLER_88_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6267_ _6234_/A _6234_/B _6266_/Y vssd1 vssd1 vccd1 vccd1 _6272_/A sky130_fd_sc_hd__a21oi_1
XFILLER_76_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8006_ _8006_/A _8006_/B vssd1 vssd1 vccd1 vccd1 _8006_/Y sky130_fd_sc_hd__nor2_1
XFILLER_57_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5218_ _4657_/A _5066_/B _5062_/X _5071_/X vssd1 vssd1 vccd1 vccd1 _5218_/X sky130_fd_sc_hd__o2bb2a_1
X_6198_ _6198_/A vssd1 vssd1 vccd1 vccd1 _6198_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5149_ _5149_/A _5149_/B _5219_/D _5149_/D vssd1 vssd1 vccd1 vccd1 _5149_/X sky130_fd_sc_hd__or4_1
XFILLER_29_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8908_ _8908_/A _4431_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[17] sky130_fd_sc_hd__ebufn_8
X_8839_ _8839_/A _4350_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[18] sky130_fd_sc_hd__ebufn_8
XFILLER_52_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4520_ _4520_/A _4520_/B _4732_/A vssd1 vssd1 vccd1 vccd1 _4542_/B sky130_fd_sc_hd__and3_1
X_4451_ _4451_/A vssd1 vssd1 vccd1 vccd1 _4456_/A sky130_fd_sc_hd__clkbuf_4
X_7170_ _7169_/A _7169_/B _7169_/C vssd1 vssd1 vccd1 vccd1 _7262_/C sky130_fd_sc_hd__a21o_1
XFILLER_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4382_ _4383_/A vssd1 vssd1 vccd1 vccd1 _4382_/Y sky130_fd_sc_hd__inv_2
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6121_ _6121_/A _6121_/B vssd1 vssd1 vccd1 vccd1 _6122_/B sky130_fd_sc_hd__nand2_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6052_ _6052_/A _6052_/B vssd1 vssd1 vccd1 vccd1 _6053_/B sky130_fd_sc_hd__nor2_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5003_ _5098_/B _5193_/C _5071_/A vssd1 vssd1 vccd1 vccd1 _5003_/X sky130_fd_sc_hd__o21a_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6954_ _7236_/B _6954_/B vssd1 vssd1 vccd1 vccd1 _7004_/A sky130_fd_sc_hd__xor2_2
XFILLER_34_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5905_ _6119_/A _5883_/A _6003_/A _6007_/A vssd1 vssd1 vccd1 vccd1 _6014_/B sky130_fd_sc_hd__o22a_1
X_6885_ _6973_/A _6885_/B vssd1 vssd1 vccd1 vccd1 _6886_/B sky130_fd_sc_hd__xnor2_1
XFILLER_14_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8624_ input3/X _8624_/D vssd1 vssd1 vccd1 vccd1 _8624_/Q sky130_fd_sc_hd__dfxtp_1
X_5836_ _5838_/B vssd1 vssd1 vccd1 vccd1 _6205_/A sky130_fd_sc_hd__clkbuf_2
X_8555_ _8556_/A _8556_/B _8556_/C vssd1 vssd1 vccd1 vccd1 _8557_/C sky130_fd_sc_hd__a21oi_1
X_5767_ _5768_/A _5768_/B _5768_/C vssd1 vssd1 vccd1 vccd1 _5856_/A sky130_fd_sc_hd__a21oi_1
X_8486_ _8486_/A _8486_/B vssd1 vssd1 vccd1 vccd1 _8487_/B sky130_fd_sc_hd__xnor2_1
X_7506_ _7508_/B _7505_/Y _7509_/A vssd1 vssd1 vccd1 vccd1 _7506_/X sky130_fd_sc_hd__o21ba_1
X_5698_ _5699_/A _5699_/B vssd1 vssd1 vccd1 vccd1 _5711_/B sky130_fd_sc_hd__nand2_1
X_4718_ _4718_/A vssd1 vssd1 vccd1 vccd1 _8599_/D sky130_fd_sc_hd__clkbuf_1
X_7437_ _7446_/A _7437_/B vssd1 vssd1 vccd1 vccd1 _7442_/A sky130_fd_sc_hd__nand2_1
X_4649_ _6507_/A vssd1 vssd1 vccd1 vccd1 _4650_/A sky130_fd_sc_hd__buf_2
X_7368_ _7368_/A _7368_/B vssd1 vssd1 vccd1 vccd1 _7395_/A sky130_fd_sc_hd__xnor2_1
X_8728__6 vssd1 vssd1 vccd1 vccd1 _8728__6/HI _8823_/A sky130_fd_sc_hd__conb_1
X_7299_ _7299_/A _7299_/B vssd1 vssd1 vccd1 vccd1 _7315_/C sky130_fd_sc_hd__xnor2_1
X_6319_ _6309_/A _6309_/B _6310_/X _6314_/Y _6318_/X vssd1 vssd1 vccd1 vccd1 _6326_/C
+ sky130_fd_sc_hd__a2111o_1
XFILLER_39_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8788__66 vssd1 vssd1 vccd1 vccd1 _8788__66/HI _8897_/A sky130_fd_sc_hd__conb_1
XFILLER_57_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6670_ _6670_/A vssd1 vssd1 vccd1 vccd1 _6700_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_31_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5621_ _8649_/Q _7634_/A vssd1 vssd1 vccd1 vccd1 _5638_/B sky130_fd_sc_hd__and2b_1
X_8340_ _8341_/A _8341_/B _8341_/C vssd1 vssd1 vccd1 vccd1 _8342_/A sky130_fd_sc_hd__a21oi_1
X_5552_ _6119_/A _5898_/A _5551_/X vssd1 vssd1 vccd1 vccd1 _5553_/B sky130_fd_sc_hd__o21a_1
X_8271_ _8255_/B _8257_/B _8255_/A vssd1 vssd1 vccd1 vccd1 _8349_/A sky130_fd_sc_hd__o21ba_1
X_4503_ _8605_/Q vssd1 vssd1 vccd1 vccd1 _7627_/B sky130_fd_sc_hd__buf_4
X_5483_ _5486_/A _5486_/B _5460_/A vssd1 vssd1 vccd1 vccd1 _5520_/B sky130_fd_sc_hd__a21oi_2
X_7222_ _6593_/A _6864_/A _7227_/A vssd1 vssd1 vccd1 vccd1 _7222_/X sky130_fd_sc_hd__o21ba_1
X_4434_ _4438_/A vssd1 vssd1 vccd1 vccd1 _4434_/Y sky130_fd_sc_hd__inv_2
X_7153_ _7153_/A _7153_/B vssd1 vssd1 vccd1 vccd1 _7155_/A sky130_fd_sc_hd__xnor2_1
X_4365_ _4365_/A vssd1 vssd1 vccd1 vccd1 _4370_/A sky130_fd_sc_hd__buf_6
X_7084_ _7084_/A _7084_/B vssd1 vssd1 vccd1 vccd1 _7147_/B sky130_fd_sc_hd__xnor2_2
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6104_ _6102_/X _6104_/B _6167_/A vssd1 vssd1 vccd1 vccd1 _6106_/A sky130_fd_sc_hd__and3b_1
XFILLER_58_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6035_ _5801_/C _6119_/A _6214_/B vssd1 vssd1 vccd1 vccd1 _6081_/B sky130_fd_sc_hd__a21bo_1
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7986_ _7986_/A _8056_/B vssd1 vssd1 vccd1 vccd1 _8166_/A sky130_fd_sc_hd__nand2_2
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6937_ _6936_/A _6936_/B _6936_/C vssd1 vssd1 vccd1 vccd1 _7044_/D sky130_fd_sc_hd__a21oi_1
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6868_ _6868_/A _6868_/B vssd1 vssd1 vccd1 vccd1 _6876_/B sky130_fd_sc_hd__xnor2_1
XFILLER_22_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5819_ _5820_/A _5820_/B _6218_/A vssd1 vssd1 vccd1 vccd1 _5875_/A sky130_fd_sc_hd__a21o_1
X_8607_ input3/X _8607_/D vssd1 vssd1 vccd1 vccd1 _8607_/Q sky130_fd_sc_hd__dfxtp_1
X_8538_ _8538_/A _8706_/Q vssd1 vssd1 vccd1 vccd1 _8540_/A sky130_fd_sc_hd__nor2_1
X_6799_ _6799_/A vssd1 vssd1 vccd1 vccd1 _7048_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_41_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8469_ _8397_/A _8397_/B _8398_/B _8194_/A vssd1 vssd1 vccd1 vccd1 _8470_/B sky130_fd_sc_hd__a22o_1
XFILLER_77_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7840_ _7887_/A _8206_/A vssd1 vssd1 vccd1 vccd1 _8508_/B sky130_fd_sc_hd__nor2_1
XFILLER_36_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7771_ _7887_/A _8331_/A _7771_/C vssd1 vssd1 vccd1 vccd1 _7772_/B sky130_fd_sc_hd__nor3_1
XFILLER_51_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4983_ _5066_/A _5092_/A _4983_/C vssd1 vssd1 vccd1 vccd1 _4983_/X sky130_fd_sc_hd__or3_1
X_6722_ _6789_/A _6722_/B vssd1 vssd1 vccd1 vccd1 _6790_/A sky130_fd_sc_hd__xnor2_1
XFILLER_51_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6653_ _6660_/A _6652_/B _6652_/C vssd1 vssd1 vccd1 vccd1 _7176_/C sky130_fd_sc_hd__a21o_1
XFILLER_31_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5604_ _5713_/A _5713_/B vssd1 vssd1 vccd1 vccd1 _6061_/A sky130_fd_sc_hd__xor2_2
X_6584_ _6592_/A _6584_/B vssd1 vssd1 vccd1 vccd1 _7193_/A sky130_fd_sc_hd__xnor2_4
X_8323_ _8381_/A _8323_/B vssd1 vssd1 vccd1 vccd1 _8343_/A sky130_fd_sc_hd__xnor2_1
X_5535_ _5800_/A _5580_/B vssd1 vssd1 vccd1 vccd1 _5560_/A sky130_fd_sc_hd__nor2_1
XFILLER_11_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8254_ _8254_/A _8254_/B _8254_/C vssd1 vssd1 vccd1 vccd1 _8255_/B sky130_fd_sc_hd__nor3_1
X_5466_ _8661_/Q _8598_/Q vssd1 vssd1 vccd1 vccd1 _5468_/A sky130_fd_sc_hd__and2b_1
X_7205_ _7205_/A _7205_/B vssd1 vssd1 vccd1 vccd1 _7206_/B sky130_fd_sc_hd__xnor2_2
X_4417_ _4420_/A vssd1 vssd1 vccd1 vccd1 _4417_/Y sky130_fd_sc_hd__inv_2
X_8185_ _8185_/A vssd1 vssd1 vccd1 vccd1 _8185_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5397_ _5414_/A _8647_/Q _5428_/A _5421_/A vssd1 vssd1 vccd1 vccd1 _5397_/X sky130_fd_sc_hd__a211o_1
X_4348_ _4352_/A vssd1 vssd1 vccd1 vccd1 _4348_/Y sky130_fd_sc_hd__inv_2
X_7136_ _7378_/B _6814_/B _7136_/S vssd1 vssd1 vccd1 vccd1 _7140_/A sky130_fd_sc_hd__mux2_1
X_7067_ _7067_/A _7135_/B vssd1 vssd1 vccd1 vccd1 _7068_/B sky130_fd_sc_hd__xnor2_1
XFILLER_74_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6018_ _6018_/A _6018_/B vssd1 vssd1 vccd1 vccd1 _6019_/B sky130_fd_sc_hd__and2_1
XFILLER_46_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8758__36 vssd1 vssd1 vccd1 vccd1 _8758__36/HI _8853_/A sky130_fd_sc_hd__conb_1
XFILLER_27_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7969_ _7969_/A _8023_/B _7969_/C vssd1 vssd1 vccd1 vccd1 _8022_/A sky130_fd_sc_hd__nand3_1
XFILLER_14_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8772__50 vssd1 vssd1 vccd1 vccd1 _8772__50/HI _8881_/A sky130_fd_sc_hd__conb_1
XFILLER_60_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5320_ _5320_/A vssd1 vssd1 vccd1 vccd1 _5354_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_5251_ _5251_/A _5251_/B vssd1 vssd1 vccd1 vccd1 _5251_/X sky130_fd_sc_hd__or2_1
X_5182_ _5194_/A _5185_/C _5182_/C vssd1 vssd1 vccd1 vccd1 _5182_/X sky130_fd_sc_hd__or3_1
XFILLER_56_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8872_ _8872_/A _4389_/Y vssd1 vssd1 vccd1 vccd1 io_out[19] sky130_fd_sc_hd__ebufn_8
XFILLER_64_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7823_ _7823_/A vssd1 vssd1 vccd1 vccd1 _8207_/A sky130_fd_sc_hd__buf_2
XFILLER_51_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7754_ _7740_/A _7740_/B _7747_/X vssd1 vssd1 vccd1 vccd1 _7766_/C sky130_fd_sc_hd__a21o_1
X_6705_ _6705_/A _6760_/A vssd1 vssd1 vccd1 vccd1 _7172_/B sky130_fd_sc_hd__xnor2_1
XFILLER_11_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4966_ _5120_/A _5241_/B vssd1 vssd1 vccd1 vccd1 _5165_/C sky130_fd_sc_hd__or2_1
X_7685_ _7685_/A _7685_/B vssd1 vssd1 vccd1 vccd1 _7685_/X sky130_fd_sc_hd__or2_1
X_4897_ _4897_/A _4897_/B _4897_/C vssd1 vssd1 vccd1 vccd1 _5159_/B sky130_fd_sc_hd__nor3_4
XFILLER_22_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6636_ _6737_/A _6737_/B _7092_/A vssd1 vssd1 vccd1 vccd1 _6772_/A sky130_fd_sc_hd__a21oi_2
X_6567_ _6567_/A _7627_/B vssd1 vssd1 vccd1 vccd1 _6591_/B sky130_fd_sc_hd__nand2_1
X_8306_ _8306_/A _8306_/B vssd1 vssd1 vccd1 vccd1 _8385_/B sky130_fd_sc_hd__nand2_1
X_5518_ _5724_/C vssd1 vssd1 vccd1 vccd1 _5794_/C sky130_fd_sc_hd__clkbuf_2
X_6498_ _8687_/Q vssd1 vssd1 vccd1 vccd1 _6526_/B sky130_fd_sc_hd__inv_2
X_8237_ _8341_/B _8237_/B vssd1 vssd1 vccd1 vccd1 _8238_/B sky130_fd_sc_hd__nand2_1
X_5449_ _5615_/A _5449_/B _5449_/C vssd1 vssd1 vccd1 vccd1 _5451_/B sky130_fd_sc_hd__or3_1
XFILLER_99_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8168_ _8371_/A _8168_/B _8168_/C vssd1 vssd1 vccd1 vccd1 _8169_/B sky130_fd_sc_hd__nand3_1
XFILLER_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7119_ _7024_/A _7024_/B _7118_/X vssd1 vssd1 vccd1 vccd1 _7120_/B sky130_fd_sc_hd__a21o_1
X_8099_ _8089_/B _8099_/B vssd1 vssd1 vccd1 vccd1 _8099_/X sky130_fd_sc_hd__and2b_1
XFILLER_74_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4820_ _4820_/A _4820_/B vssd1 vssd1 vccd1 vccd1 _4836_/B sky130_fd_sc_hd__nand2_4
XFILLER_33_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4751_ _4824_/C _4897_/A vssd1 vssd1 vccd1 vccd1 _4752_/A sky130_fd_sc_hd__or2_1
X_7470_ _7470_/A _7470_/B vssd1 vssd1 vccd1 vccd1 _7508_/A sky130_fd_sc_hd__xnor2_2
X_4682_ _4710_/A vssd1 vssd1 vccd1 vccd1 _4707_/A sky130_fd_sc_hd__clkbuf_1
X_6421_ _6397_/D _6422_/C _6420_/Y vssd1 vssd1 vccd1 vccd1 _8669_/D sky130_fd_sc_hd__a21oi_1
X_6352_ _6352_/A _6352_/B vssd1 vssd1 vccd1 vccd1 _6354_/A sky130_fd_sc_hd__nor2_1
X_5303_ _8628_/Q vssd1 vssd1 vccd1 vccd1 _6475_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6283_ _5754_/B _5985_/A _6204_/B _5956_/B vssd1 vssd1 vccd1 vccd1 _6285_/A sky130_fd_sc_hd__a211o_1
XFILLER_102_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8022_ _8022_/A _8022_/B vssd1 vssd1 vccd1 vccd1 _8105_/B sky130_fd_sc_hd__nand2_1
XFILLER_69_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5234_ _5234_/A _5253_/B _5234_/C vssd1 vssd1 vccd1 vccd1 _5234_/X sky130_fd_sc_hd__or3_1
X_5165_ _5219_/A _5219_/B _5165_/C _5165_/D vssd1 vssd1 vccd1 vccd1 _5165_/X sky130_fd_sc_hd__or4_1
XFILLER_83_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5096_ _5215_/D _5096_/B vssd1 vssd1 vccd1 vccd1 _5096_/X sky130_fd_sc_hd__or2_1
XFILLER_29_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8924_ _8924_/A _4450_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[33] sky130_fd_sc_hd__ebufn_8
XFILLER_56_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8855_ _8855_/A _4368_/Y vssd1 vssd1 vccd1 vccd1 io_out[2] sky130_fd_sc_hd__ebufn_8
XFILLER_71_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7806_ _7807_/A _7807_/B vssd1 vssd1 vccd1 vccd1 _7851_/A sky130_fd_sc_hd__nor2_1
XFILLER_52_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5998_ _5998_/A _6202_/A vssd1 vssd1 vccd1 vccd1 _6000_/B sky130_fd_sc_hd__xnor2_1
X_7737_ _7869_/A _7869_/B vssd1 vssd1 vccd1 vccd1 _7864_/B sky130_fd_sc_hd__xor2_1
X_4949_ _4657_/A _5135_/C _5176_/B _4948_/X vssd1 vssd1 vccd1 vccd1 _4949_/X sky130_fd_sc_hd__o31a_1
XFILLER_24_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7668_ _7816_/A _7668_/B vssd1 vssd1 vccd1 vccd1 _7819_/B sky130_fd_sc_hd__xnor2_1
X_6619_ _8691_/Q _8608_/Q vssd1 vssd1 vccd1 vccd1 _6660_/B sky130_fd_sc_hd__or2b_1
XFILLER_20_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7599_ _7599_/A vssd1 vssd1 vccd1 vccd1 _8710_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8742__20 vssd1 vssd1 vccd1 vccd1 _8742__20/HI _8837_/A sky130_fd_sc_hd__conb_1
XFILLER_30_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6970_ _6850_/A _6970_/B vssd1 vssd1 vccd1 vccd1 _6970_/X sky130_fd_sc_hd__and2b_1
X_5921_ _6193_/A _5921_/B vssd1 vssd1 vccd1 vccd1 _5950_/A sky130_fd_sc_hd__nand2_1
XFILLER_19_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5852_ _5850_/Y _5852_/B vssd1 vssd1 vccd1 vccd1 _5937_/B sky130_fd_sc_hd__and2b_1
XFILLER_34_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8640_ input3/X _8640_/D vssd1 vssd1 vccd1 vccd1 _8640_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4803_ _4820_/A _4803_/B _4872_/A vssd1 vssd1 vccd1 vccd1 _4829_/A sky130_fd_sc_hd__or3_1
X_5783_ _5783_/A _5861_/B vssd1 vssd1 vccd1 vccd1 _6032_/B sky130_fd_sc_hd__xnor2_1
X_8571_ input3/X _8571_/D vssd1 vssd1 vccd1 vccd1 _8571_/Q sky130_fd_sc_hd__dfxtp_1
X_7522_ _7522_/A _7522_/B vssd1 vssd1 vccd1 vccd1 _7522_/X sky130_fd_sc_hd__xor2_1
X_4734_ _6406_/A vssd1 vssd1 vccd1 vccd1 _7503_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_9_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7453_ _7482_/A _7482_/B _7478_/A _7477_/A vssd1 vssd1 vccd1 vccd1 _7480_/C sky130_fd_sc_hd__o211ai_2
X_4665_ _8593_/Q vssd1 vssd1 vccd1 vccd1 _5068_/A sky130_fd_sc_hd__inv_2
X_7384_ _7385_/A _7385_/B vssd1 vssd1 vccd1 vccd1 _7384_/Y sky130_fd_sc_hd__nor2_1
X_4596_ _8574_/Q _4598_/C _4595_/X vssd1 vssd1 vccd1 vccd1 _4597_/B sky130_fd_sc_hd__o21ai_1
X_6404_ _8665_/Q _6468_/B vssd1 vssd1 vccd1 vccd1 _6405_/A sky130_fd_sc_hd__and2b_1
X_6335_ _6329_/X _6333_/X _6334_/X _8655_/Q vssd1 vssd1 vccd1 vccd1 _8655_/D sky130_fd_sc_hd__o2bb2a_1
X_8005_ _8006_/A _8006_/B vssd1 vssd1 vccd1 vccd1 _8083_/A sky130_fd_sc_hd__and2_1
X_6266_ _6266_/A _6266_/B vssd1 vssd1 vccd1 vccd1 _6266_/Y sky130_fd_sc_hd__nor2_1
XFILLER_88_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6197_ _6197_/A _6197_/B vssd1 vssd1 vccd1 vccd1 _6239_/A sky130_fd_sc_hd__xnor2_2
X_5217_ _5053_/D _5070_/D _5072_/X _5216_/X vssd1 vssd1 vccd1 vccd1 _5217_/X sky130_fd_sc_hd__o31a_1
XFILLER_96_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5148_ _5251_/A _5136_/X _5140_/X _5190_/A _5147_/Y vssd1 vssd1 vccd1 vccd1 _5148_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_17_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5079_ _5143_/A _5224_/D vssd1 vssd1 vccd1 vccd1 _5079_/X sky130_fd_sc_hd__and2_1
XFILLER_84_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8907_ _8907_/A _4430_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[16] sky130_fd_sc_hd__ebufn_8
XFILLER_44_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8838_ _8838_/A _4349_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[17] sky130_fd_sc_hd__ebufn_8
XFILLER_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4450_ _4450_/A vssd1 vssd1 vccd1 vccd1 _4450_/Y sky130_fd_sc_hd__inv_2
X_4381_ _4383_/A vssd1 vssd1 vccd1 vccd1 _4381_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6120_ _6121_/A _6121_/B vssd1 vssd1 vccd1 vccd1 _6135_/B sky130_fd_sc_hd__or2_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6051_ _6050_/B _6051_/B vssd1 vssd1 vccd1 vccd1 _6052_/B sky130_fd_sc_hd__and2b_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5002_ _5102_/C _5122_/B vssd1 vssd1 vccd1 vccd1 _5193_/C sky130_fd_sc_hd__or2_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6953_ _7039_/A _7039_/B vssd1 vssd1 vccd1 vccd1 _6961_/A sky130_fd_sc_hd__xnor2_1
XFILLER_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6884_ _7006_/A _6884_/B vssd1 vssd1 vccd1 vccd1 _6885_/B sky130_fd_sc_hd__xnor2_1
XFILLER_81_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5904_ _5812_/A _6220_/B _5805_/A _5903_/A vssd1 vssd1 vccd1 vccd1 _5912_/B sky130_fd_sc_hd__o211ai_1
X_8623_ input3/X _8623_/D vssd1 vssd1 vccd1 vccd1 _8623_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5835_ _5954_/A _5954_/C _5956_/B vssd1 vssd1 vccd1 vccd1 _5838_/B sky130_fd_sc_hd__o21ba_1
XFILLER_22_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8554_ _7702_/Y _8561_/B _8553_/X vssd1 vssd1 vccd1 vccd1 _8556_/C sky130_fd_sc_hd__a21oi_1
X_5766_ _5824_/A _5824_/B vssd1 vssd1 vccd1 vccd1 _5768_/C sky130_fd_sc_hd__xnor2_1
X_8485_ _8485_/A _8485_/B vssd1 vssd1 vccd1 vccd1 _8486_/B sky130_fd_sc_hd__xnor2_1
X_7505_ _7505_/A _7505_/B _7505_/C vssd1 vssd1 vccd1 vccd1 _7505_/Y sky130_fd_sc_hd__nor3_1
X_5697_ _5697_/A _5697_/B vssd1 vssd1 vccd1 vccd1 _5699_/B sky130_fd_sc_hd__xnor2_1
X_4717_ _4717_/A _4717_/B _4724_/S vssd1 vssd1 vccd1 vccd1 _4718_/A sky130_fd_sc_hd__and3_1
X_7436_ _7436_/A _7436_/B vssd1 vssd1 vccd1 vccd1 _7437_/B sky130_fd_sc_hd__or2_1
XFILLER_30_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4648_ _4648_/A vssd1 vssd1 vccd1 vccd1 _6507_/A sky130_fd_sc_hd__clkbuf_4
X_7367_ _7367_/A _7367_/B vssd1 vssd1 vccd1 vccd1 _7480_/A sky130_fd_sc_hd__nor2_1
XFILLER_1_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4579_ _8579_/Q _4579_/B _4579_/C vssd1 vssd1 vccd1 vccd1 _5406_/B sky130_fd_sc_hd__or3_4
X_7298_ _7315_/A _7314_/A vssd1 vssd1 vccd1 vccd1 _7300_/A sky130_fd_sc_hd__nand2_1
XFILLER_1_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6318_ _6314_/A _6314_/B _6315_/X _6316_/Y _6317_/X vssd1 vssd1 vccd1 vccd1 _6318_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_103_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6249_ _6249_/A _6249_/B vssd1 vssd1 vccd1 vccd1 _6249_/Y sky130_fd_sc_hd__nand2_1
XFILLER_39_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5620_ _5620_/A _8649_/Q vssd1 vssd1 vccd1 vccd1 _5680_/A sky130_fd_sc_hd__or2b_1
XFILLER_31_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5551_ _5551_/A _6003_/A vssd1 vssd1 vccd1 vccd1 _5551_/X sky130_fd_sc_hd__or2_1
X_8270_ _8260_/A _8260_/B _8269_/Y vssd1 vssd1 vccd1 vccd1 _8429_/A sky130_fd_sc_hd__a21o_1
XFILLER_8_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4502_ _4802_/B _4842_/C vssd1 vssd1 vccd1 vccd1 _4822_/A sky130_fd_sc_hd__and2_1
X_7221_ _7223_/B _7289_/B vssd1 vssd1 vccd1 vccd1 _7230_/A sky130_fd_sc_hd__xor2_1
X_5482_ _5482_/A _5482_/B vssd1 vssd1 vccd1 vccd1 _5520_/A sky130_fd_sc_hd__nand2_2
X_4433_ _4451_/A vssd1 vssd1 vccd1 vccd1 _4438_/A sky130_fd_sc_hd__buf_2
XFILLER_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4364_ _4364_/A vssd1 vssd1 vccd1 vccd1 _4364_/Y sky130_fd_sc_hd__inv_2
X_7152_ _7008_/A _7006_/X _7030_/B _6880_/A vssd1 vssd1 vccd1 vccd1 _7153_/B sky130_fd_sc_hd__a2bb2o_1
X_7083_ _7083_/A _7083_/B vssd1 vssd1 vccd1 vccd1 _7084_/B sky130_fd_sc_hd__nor2_1
XFILLER_86_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6103_ _6103_/A _6103_/B _6103_/C vssd1 vssd1 vccd1 vccd1 _6104_/B sky130_fd_sc_hd__or3_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6034_ _6034_/A _6034_/B vssd1 vssd1 vccd1 vccd1 _6214_/B sky130_fd_sc_hd__and2_1
XFILLER_100_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7985_ _8051_/A _8384_/A _7985_/C vssd1 vssd1 vccd1 vccd1 _7992_/B sky130_fd_sc_hd__and3_1
XFILLER_26_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6936_ _6936_/A _6936_/B _6936_/C vssd1 vssd1 vccd1 vccd1 _7044_/C sky130_fd_sc_hd__and3_1
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6867_ _6880_/A _6880_/B vssd1 vssd1 vccd1 vccd1 _6868_/B sky130_fd_sc_hd__xnor2_1
XFILLER_34_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8730__8 vssd1 vssd1 vccd1 vccd1 _8730__8/HI _8825_/A sky130_fd_sc_hd__conb_1
X_6798_ _6798_/A _6798_/B vssd1 vssd1 vccd1 vccd1 _7060_/A sky130_fd_sc_hd__nor2_2
X_5818_ _5997_/A _5803_/B _6259_/A vssd1 vssd1 vccd1 vccd1 _6218_/A sky130_fd_sc_hd__o21ai_4
X_8606_ input3/X _8606_/D vssd1 vssd1 vccd1 vccd1 _8606_/Q sky130_fd_sc_hd__dfxtp_4
X_8537_ _8537_/A vssd1 vssd1 vccd1 vccd1 _8720_/D sky130_fd_sc_hd__clkbuf_1
X_5749_ _5754_/A _5749_/B vssd1 vssd1 vccd1 vccd1 _5849_/B sky130_fd_sc_hd__nand2_1
X_8468_ _8407_/S _8408_/A _8467_/X vssd1 vssd1 vccd1 vccd1 _8470_/A sky130_fd_sc_hd__a21bo_1
X_8399_ _8400_/A _8400_/B _8400_/C vssd1 vssd1 vccd1 vccd1 _8401_/A sky130_fd_sc_hd__o21ai_1
X_7419_ _7418_/A _7418_/B _7418_/C vssd1 vssd1 vccd1 vccd1 _7420_/B sky130_fd_sc_hd__a21oi_1
XFILLER_104_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7770_ _8205_/B _8327_/A vssd1 vssd1 vccd1 vccd1 _7771_/C sky130_fd_sc_hd__nor2_1
X_4982_ _5091_/D _4977_/X _4981_/X _4657_/A vssd1 vssd1 vccd1 vccd1 _4983_/C sky130_fd_sc_hd__o22a_1
X_6721_ _6951_/A _6805_/A vssd1 vssd1 vccd1 vccd1 _6722_/B sky130_fd_sc_hd__xnor2_1
XFILLER_23_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6652_ _6660_/A _6652_/B _6652_/C vssd1 vssd1 vccd1 vccd1 _7176_/B sky130_fd_sc_hd__nand3_1
X_5603_ _5603_/A _5603_/B vssd1 vssd1 vccd1 vccd1 _5713_/B sky130_fd_sc_hd__xor2_2
X_8322_ _8322_/A _8380_/A vssd1 vssd1 vccd1 vccd1 _8323_/B sky130_fd_sc_hd__xnor2_1
X_6583_ _7175_/A _7238_/A vssd1 vssd1 vccd1 vccd1 _6815_/B sky130_fd_sc_hd__nand2_1
XFILLER_11_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5534_ _5584_/A _5534_/B vssd1 vssd1 vccd1 vccd1 _5800_/A sky130_fd_sc_hd__xnor2_4
X_8253_ _8254_/A _8254_/B _8254_/C vssd1 vssd1 vccd1 vccd1 _8255_/A sky130_fd_sc_hd__o21a_1
X_5465_ _5584_/A _5534_/B _5464_/X vssd1 vssd1 vccd1 vccd1 _5475_/B sky130_fd_sc_hd__a21o_1
X_7204_ _7187_/A _7187_/B _7203_/X vssd1 vssd1 vccd1 vccd1 _7206_/A sky130_fd_sc_hd__a21bo_1
X_8184_ _8264_/A _8264_/B vssd1 vssd1 vccd1 vccd1 _8262_/A sky130_fd_sc_hd__and2_1
X_4416_ _4420_/A vssd1 vssd1 vccd1 vccd1 _4416_/Y sky130_fd_sc_hd__inv_2
X_7135_ _7135_/A _7135_/B vssd1 vssd1 vccd1 vccd1 _7136_/S sky130_fd_sc_hd__nand2_1
X_5396_ _8649_/Q vssd1 vssd1 vccd1 vccd1 _5421_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_101_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4347_ _4365_/A vssd1 vssd1 vccd1 vccd1 _4352_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_86_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7066_ _7239_/A _7114_/B vssd1 vssd1 vccd1 vccd1 _7135_/B sky130_fd_sc_hd__xnor2_1
XFILLER_59_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6017_ _6231_/A _6017_/B _6231_/B vssd1 vssd1 vccd1 vccd1 _6018_/B sky130_fd_sc_hd__nand3_1
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7968_ _8023_/A _7967_/B _7967_/C vssd1 vssd1 vccd1 vccd1 _7969_/C sky130_fd_sc_hd__a21o_1
XFILLER_27_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7899_ _8207_/A _8331_/A _7898_/C _7898_/D vssd1 vssd1 vccd1 vccd1 _7948_/C sky130_fd_sc_hd__a22o_1
X_6919_ _6919_/A _6919_/B _7177_/A vssd1 vssd1 vccd1 vccd1 _7062_/A sky130_fd_sc_hd__or3_1
XFILLER_52_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5250_ _4728_/B _5109_/B _5244_/X _5249_/X _4728_/A vssd1 vssd1 vccd1 vccd1 _5251_/B
+ sky130_fd_sc_hd__o32a_1
XFILLER_87_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5181_ _5183_/S _5185_/C _5132_/B _5118_/D _5180_/X vssd1 vssd1 vccd1 vccd1 _5181_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8871_ _8871_/A _4388_/Y vssd1 vssd1 vccd1 vccd1 io_out[18] sky130_fd_sc_hd__ebufn_8
XFILLER_91_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7822_ _7833_/A _7822_/B vssd1 vssd1 vccd1 vccd1 _7841_/A sky130_fd_sc_hd__nand2_1
XFILLER_64_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7753_ _7753_/A _8561_/A vssd1 vssd1 vccd1 vccd1 _7766_/A sky130_fd_sc_hd__or2b_2
XFILLER_51_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4965_ _5145_/B _5076_/A vssd1 vssd1 vccd1 vccd1 _5086_/A sky130_fd_sc_hd__or2_1
X_6704_ _7163_/B _7163_/C _7163_/A vssd1 vssd1 vccd1 vccd1 _6760_/A sky130_fd_sc_hd__a21boi_2
X_7684_ _7904_/A _8301_/A _7683_/C vssd1 vssd1 vccd1 vccd1 _7685_/B sky130_fd_sc_hd__a21oi_1
X_4896_ _5193_/B vssd1 vssd1 vccd1 vccd1 _5151_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6635_ _6635_/A vssd1 vssd1 vccd1 vccd1 _7092_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6566_ _6566_/A vssd1 vssd1 vccd1 vccd1 _6591_/A sky130_fd_sc_hd__buf_2
X_8305_ _8305_/A _8305_/B vssd1 vssd1 vccd1 vccd1 _8384_/B sky130_fd_sc_hd__or2_1
XFILLER_3_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5517_ _5724_/B vssd1 vssd1 vccd1 vccd1 _5794_/B sky130_fd_sc_hd__clkbuf_2
X_8236_ _8236_/A _8236_/B vssd1 vssd1 vccd1 vccd1 _8237_/B sky130_fd_sc_hd__nand2_1
X_6497_ _6520_/A _6514_/A _6526_/A vssd1 vssd1 vccd1 vccd1 _6497_/X sky130_fd_sc_hd__o21a_1
X_5448_ _5447_/X _5442_/C _5448_/S vssd1 vssd1 vccd1 vccd1 _5449_/C sky130_fd_sc_hd__mux2_1
X_8818__96 vssd1 vssd1 vccd1 vccd1 _8818__96/HI _8927_/A sky130_fd_sc_hd__conb_1
XFILLER_87_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8167_ _8168_/B _8168_/C _8371_/A vssd1 vssd1 vccd1 vccd1 _8293_/A sky130_fd_sc_hd__a21o_1
XFILLER_59_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5379_ _8660_/Q vssd1 vssd1 vccd1 vccd1 _5462_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_7118_ _7131_/A _7118_/B vssd1 vssd1 vccd1 vccd1 _7118_/X sky130_fd_sc_hd__and2_1
X_8098_ _8499_/A _8501_/A _8499_/B vssd1 vssd1 vccd1 vccd1 _8503_/C sky130_fd_sc_hd__a21o_1
XFILLER_59_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7049_ _7045_/B _6905_/B _7048_/X vssd1 vssd1 vccd1 vccd1 _7049_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_86_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4750_ _4787_/B vssd1 vssd1 vccd1 vccd1 _4897_/A sky130_fd_sc_hd__clkbuf_2
X_4681_ _4739_/A _4681_/B vssd1 vssd1 vccd1 vccd1 _4710_/A sky130_fd_sc_hd__nand2_1
X_6420_ _6397_/D _6422_/C _6419_/X vssd1 vssd1 vccd1 vccd1 _6420_/Y sky130_fd_sc_hd__o21ai_1
X_6351_ _6351_/A _8645_/Q vssd1 vssd1 vccd1 vccd1 _6352_/B sky130_fd_sc_hd__and2_1
X_5302_ _8625_/Q _8624_/Q vssd1 vssd1 vccd1 vccd1 _6478_/A sky130_fd_sc_hd__or2_1
X_6282_ _6187_/A _6187_/B _6281_/X vssd1 vssd1 vccd1 vccd1 _6286_/A sky130_fd_sc_hd__a21oi_1
XFILLER_102_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8021_ _8021_/A _8021_/B vssd1 vssd1 vccd1 vccd1 _8103_/A sky130_fd_sc_hd__nand2_1
X_5233_ _5077_/Y _5230_/X _5231_/X _5232_/X vssd1 vssd1 vccd1 vccd1 _5234_/C sky130_fd_sc_hd__o2bb2a_1
X_5164_ _4990_/A _5151_/B _5173_/B _5046_/B _5163_/Y vssd1 vssd1 vccd1 vccd1 _5165_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_68_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5095_ _5215_/B _5166_/D _5012_/A _5094_/X _4916_/B vssd1 vssd1 vccd1 vccd1 _5096_/B
+ sky130_fd_sc_hd__o32a_1
X_8923_ _8923_/A _4449_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[32] sky130_fd_sc_hd__ebufn_8
XFILLER_83_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8854_ _8854_/A _4367_/Y vssd1 vssd1 vccd1 vccd1 io_out[1] sky130_fd_sc_hd__ebufn_8
XFILLER_83_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7805_ _7936_/A _7805_/B vssd1 vssd1 vccd1 vccd1 _7807_/B sky130_fd_sc_hd__nand2_1
XFILLER_64_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5997_ _5997_/A _5997_/B vssd1 vssd1 vccd1 vccd1 _6202_/A sky130_fd_sc_hd__xnor2_1
X_7736_ _7740_/A _7740_/B _7747_/A vssd1 vssd1 vccd1 vccd1 _7869_/B sky130_fd_sc_hd__a21oi_2
X_4948_ _5183_/S _5202_/A _5202_/B _5173_/B vssd1 vssd1 vccd1 vccd1 _4948_/X sky130_fd_sc_hd__or4_1
X_7667_ _7651_/Y _7819_/A _7666_/X vssd1 vssd1 vccd1 vccd1 _7668_/B sky130_fd_sc_hd__a21oi_1
X_4879_ _5023_/A _5193_/B vssd1 vssd1 vccd1 vccd1 _5130_/B sky130_fd_sc_hd__or2_1
X_6618_ _8690_/Q _7634_/A vssd1 vssd1 vccd1 vccd1 _6620_/A sky130_fd_sc_hd__or2b_1
XFILLER_20_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7598_ _8536_/A _7598_/B vssd1 vssd1 vccd1 vccd1 _7599_/A sky130_fd_sc_hd__and2_1
XFILLER_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6549_ _7547_/A _6549_/B _6549_/C vssd1 vssd1 vccd1 vccd1 _6550_/A sky130_fd_sc_hd__and3_1
X_8219_ _8127_/A _8127_/B _8218_/X vssd1 vssd1 vccd1 vccd1 _8224_/A sky130_fd_sc_hd__a21oi_1
XFILLER_87_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5920_ _5920_/A _5920_/B _5920_/C vssd1 vssd1 vccd1 vccd1 _5935_/A sky130_fd_sc_hd__and3_1
XFILLER_34_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5851_ _5850_/A _5850_/C _5850_/B vssd1 vssd1 vccd1 vccd1 _5852_/B sky130_fd_sc_hd__o21ai_1
X_8570_ _7875_/A _8568_/Y _8569_/Y vssd1 vssd1 vccd1 vccd1 _8725_/D sky130_fd_sc_hd__a21oi_1
X_4802_ _4824_/B _4802_/B _4909_/A _4831_/A vssd1 vssd1 vccd1 vccd1 _4860_/A sky130_fd_sc_hd__or4b_2
X_5782_ _5858_/A _5782_/B vssd1 vssd1 vccd1 vccd1 _5861_/B sky130_fd_sc_hd__nand2_1
X_7521_ _7511_/S _7516_/B _7515_/A vssd1 vssd1 vccd1 vccd1 _7522_/B sky130_fd_sc_hd__o21ai_1
X_4733_ _4909_/A _4739_/B vssd1 vssd1 vccd1 vccd1 _4733_/Y sky130_fd_sc_hd__nor2_1
X_7452_ _7452_/A _7452_/B vssd1 vssd1 vccd1 vccd1 _7477_/A sky130_fd_sc_hd__or2_1
X_4664_ _4699_/B vssd1 vssd1 vccd1 vccd1 _5113_/A sky130_fd_sc_hd__clkbuf_2
X_6403_ _6419_/A vssd1 vssd1 vccd1 vccd1 _6468_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_7383_ _7374_/X _7381_/Y _7382_/X _7333_/Y vssd1 vssd1 vccd1 vccd1 _7388_/A sky130_fd_sc_hd__a211oi_1
X_4595_ _4639_/B vssd1 vssd1 vccd1 vccd1 _4595_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6334_ _7503_/A vssd1 vssd1 vccd1 vccd1 _6334_/X sky130_fd_sc_hd__buf_2
XFILLER_103_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6265_ _5828_/A _6203_/B _6204_/A vssd1 vssd1 vccd1 vccd1 _6273_/A sky130_fd_sc_hd__a21oi_1
XFILLER_103_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8004_ _8020_/B _8002_/Y _7948_/X _7929_/X vssd1 vssd1 vccd1 vccd1 _8009_/B sky130_fd_sc_hd__a211o_1
X_5216_ _5166_/D _5091_/X _5214_/X _5215_/X vssd1 vssd1 vccd1 vccd1 _5216_/X sky130_fd_sc_hd__o211a_1
X_6196_ _6196_/A vssd1 vssd1 vccd1 vccd1 _6197_/B sky130_fd_sc_hd__inv_2
XFILLER_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5147_ _5251_/A _5147_/B vssd1 vssd1 vccd1 vccd1 _5147_/Y sky130_fd_sc_hd__nand2_1
XFILLER_56_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5078_ _5017_/B _5077_/Y _5054_/C _5115_/B vssd1 vssd1 vccd1 vccd1 _5224_/D sky130_fd_sc_hd__a211o_1
X_8906_ _8906_/A _4429_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[15] sky130_fd_sc_hd__ebufn_8
XFILLER_56_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8837_ _8837_/A _4348_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[16] sky130_fd_sc_hd__ebufn_8
XFILLER_71_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7719_ _7957_/A vssd1 vssd1 vccd1 vccd1 _8116_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_12_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8699_ input3/X _8699_/D vssd1 vssd1 vccd1 vccd1 _8699_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_60_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8802__80 vssd1 vssd1 vccd1 vccd1 _8802__80/HI _8911_/A sky130_fd_sc_hd__conb_1
XFILLER_35_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4380_ _4383_/A vssd1 vssd1 vccd1 vccd1 _4380_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6050_ _6051_/B _6050_/B vssd1 vssd1 vccd1 vccd1 _6052_/A sky130_fd_sc_hd__and2b_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5001_ _4914_/X _4954_/X _5000_/X vssd1 vssd1 vccd1 vccd1 _5001_/X sky130_fd_sc_hd__a21o_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6952_ _6833_/A _6833_/B _6951_/X vssd1 vssd1 vccd1 vccd1 _7039_/B sky130_fd_sc_hd__a21oi_2
XFILLER_19_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6883_ _6947_/B _6883_/B vssd1 vssd1 vccd1 vccd1 _6884_/B sky130_fd_sc_hd__xor2_2
X_5903_ _5903_/A vssd1 vssd1 vccd1 vccd1 _6231_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_8622_ input3/X _8622_/D vssd1 vssd1 vccd1 vccd1 _8622_/Q sky130_fd_sc_hd__dfxtp_1
X_5834_ _5962_/A vssd1 vssd1 vccd1 vccd1 _5956_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_22_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8553_ _7702_/Y _8561_/B _8547_/Y vssd1 vssd1 vccd1 vccd1 _8553_/X sky130_fd_sc_hd__o21a_1
X_5765_ _5675_/A _5675_/B _5764_/X vssd1 vssd1 vccd1 vccd1 _5824_/B sky130_fd_sc_hd__a21oi_1
X_8484_ _7666_/A _8445_/A _8363_/B _8281_/Y _8147_/A vssd1 vssd1 vccd1 vccd1 _8485_/B
+ sky130_fd_sc_hd__a32o_1
X_7504_ _7505_/A _7505_/C _7505_/B vssd1 vssd1 vccd1 vccd1 _7508_/B sky130_fd_sc_hd__o21a_1
X_5696_ _6051_/B _6041_/B vssd1 vssd1 vccd1 vccd1 _5699_/A sky130_fd_sc_hd__nor2_1
X_4716_ _5226_/A _4716_/B vssd1 vssd1 vccd1 vccd1 _4724_/S sky130_fd_sc_hd__nand2_1
X_7435_ _7436_/A _7436_/B vssd1 vssd1 vccd1 vccd1 _7446_/A sky130_fd_sc_hd__nand2_1
XFILLER_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4647_ _4647_/A vssd1 vssd1 vccd1 vccd1 _8590_/D sky130_fd_sc_hd__clkbuf_1
X_7366_ _7366_/A _7366_/B _7366_/C vssd1 vssd1 vccd1 vccd1 _7367_/B sky130_fd_sc_hd__and3_1
XFILLER_89_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4578_ _4587_/A _4578_/B _4578_/C _4578_/D vssd1 vssd1 vccd1 vccd1 _4579_/C sky130_fd_sc_hd__or4_1
X_6317_ _6317_/A _6317_/B vssd1 vssd1 vccd1 vccd1 _6317_/X sky130_fd_sc_hd__xor2_2
X_7297_ _7297_/A _7297_/B vssd1 vssd1 vccd1 vccd1 _7314_/A sky130_fd_sc_hd__nor2_1
X_6248_ _6269_/A _6201_/B _6209_/B _6208_/A vssd1 vssd1 vccd1 vccd1 _6264_/A sky130_fd_sc_hd__o31a_1
X_6179_ _5967_/A _5967_/B _6178_/X vssd1 vssd1 vccd1 vccd1 _6189_/A sky130_fd_sc_hd__a21o_1
XFILLER_84_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8779__57 vssd1 vssd1 vccd1 vccd1 _8779__57/HI _8888_/A sky130_fd_sc_hd__conb_1
XFILLER_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5550_ _5507_/A _5506_/B _5507_/B _5499_/A _5549_/Y vssd1 vssd1 vccd1 vccd1 _6003_/A
+ sky130_fd_sc_hd__o311a_2
X_4501_ _8602_/Q vssd1 vssd1 vccd1 vccd1 _4842_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_5481_ _8663_/Q _8600_/Q vssd1 vssd1 vccd1 vccd1 _5482_/B sky130_fd_sc_hd__or2b_1
X_7220_ _7220_/A _7220_/B vssd1 vssd1 vccd1 vccd1 _7341_/A sky130_fd_sc_hd__xnor2_2
X_4432_ _4432_/A vssd1 vssd1 vccd1 vccd1 _4432_/Y sky130_fd_sc_hd__inv_2
XFILLER_104_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7151_ _7151_/A _7151_/B vssd1 vssd1 vccd1 vccd1 _7153_/A sky130_fd_sc_hd__xnor2_1
X_4363_ _4364_/A vssd1 vssd1 vccd1 vccd1 _4363_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7082_ _7081_/A _7081_/B _7081_/C vssd1 vssd1 vccd1 vccd1 _7083_/B sky130_fd_sc_hd__o21a_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6102_ _6161_/A _6161_/B vssd1 vssd1 vccd1 vccd1 _6102_/X sky130_fd_sc_hd__or2b_1
XFILLER_100_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6033_ _6033_/A _6033_/B vssd1 vssd1 vccd1 vccd1 _6081_/A sky130_fd_sc_hd__xnor2_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7984_ _7916_/A _7984_/B vssd1 vssd1 vccd1 vccd1 _8068_/A sky130_fd_sc_hd__and2b_1
XFILLER_26_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6935_ _6950_/A _6812_/B _6934_/X vssd1 vssd1 vccd1 vccd1 _6936_/C sky130_fd_sc_hd__a21o_1
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8793__71 vssd1 vssd1 vccd1 vccd1 _8793__71/HI _8902_/A sky130_fd_sc_hd__conb_1
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6866_ _7006_/A _6866_/B vssd1 vssd1 vccd1 vccd1 _6880_/B sky130_fd_sc_hd__xnor2_1
XFILLER_22_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6797_ _7060_/B _7099_/A vssd1 vssd1 vccd1 vccd1 _6803_/A sky130_fd_sc_hd__nor2_1
X_8605_ input3/X _8605_/D vssd1 vssd1 vccd1 vccd1 _8605_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_10_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5817_ _6323_/A _5895_/A vssd1 vssd1 vccd1 vccd1 _6259_/A sky130_fd_sc_hd__nand2_2
X_5748_ _5984_/A vssd1 vssd1 vccd1 vccd1 _6180_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_22_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8536_ _8536_/A _8536_/B vssd1 vssd1 vccd1 vccd1 _8537_/A sky130_fd_sc_hd__and2_1
X_8467_ _8395_/A _8031_/A _8407_/S _8408_/A _8408_/B vssd1 vssd1 vccd1 vccd1 _8467_/X
+ sky130_fd_sc_hd__a32o_1
X_5679_ _5679_/A _5679_/B vssd1 vssd1 vccd1 vccd1 _5680_/C sky130_fd_sc_hd__nand2_1
X_8398_ _8398_/A _8398_/B vssd1 vssd1 vccd1 vccd1 _8400_/C sky130_fd_sc_hd__xnor2_1
X_7418_ _7418_/A _7418_/B _7418_/C vssd1 vssd1 vccd1 vccd1 _7420_/A sky130_fd_sc_hd__and3_1
X_7349_ _7390_/A _7390_/B _7348_/A vssd1 vssd1 vccd1 vccd1 _7357_/A sky130_fd_sc_hd__o21bai_1
XFILLER_103_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4981_ _5098_/B _5132_/B _5055_/B _4981_/D vssd1 vssd1 vccd1 vccd1 _4981_/X sky130_fd_sc_hd__or4_1
XFILLER_23_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6720_ _7060_/B _6900_/A vssd1 vssd1 vccd1 vccd1 _6805_/A sky130_fd_sc_hd__xnor2_2
XFILLER_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6651_ _7161_/A _6651_/B vssd1 vssd1 vccd1 vccd1 _7172_/A sky130_fd_sc_hd__xnor2_1
XFILLER_31_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6582_ _6671_/A vssd1 vssd1 vccd1 vccd1 _7238_/A sky130_fd_sc_hd__clkbuf_2
X_5602_ _5602_/A _5715_/B vssd1 vssd1 vccd1 vccd1 _5603_/B sky130_fd_sc_hd__xnor2_2
X_8321_ _8321_/A _8321_/B vssd1 vssd1 vccd1 vccd1 _8380_/A sky130_fd_sc_hd__xnor2_1
X_5533_ _5539_/A _5533_/B vssd1 vssd1 vccd1 vccd1 _5551_/A sky130_fd_sc_hd__nor2_2
X_8252_ _8298_/A _8252_/B vssd1 vssd1 vccd1 vccd1 _8254_/C sky130_fd_sc_hd__and2b_1
X_5464_ _8659_/Q _8596_/Q vssd1 vssd1 vccd1 vccd1 _5464_/X sky130_fd_sc_hd__and2b_1
X_7203_ _7262_/B _7186_/B vssd1 vssd1 vccd1 vccd1 _7203_/X sky130_fd_sc_hd__or2b_1
X_8183_ _8185_/A _8183_/B vssd1 vssd1 vccd1 vccd1 _8264_/B sky130_fd_sc_hd__xnor2_1
X_4415_ _4427_/A vssd1 vssd1 vccd1 vccd1 _4420_/A sky130_fd_sc_hd__buf_2
X_5395_ _8650_/Q vssd1 vssd1 vccd1 vccd1 _5428_/A sky130_fd_sc_hd__clkbuf_2
X_4346_ _4346_/A vssd1 vssd1 vccd1 vccd1 _4346_/Y sky130_fd_sc_hd__inv_2
X_7134_ _7115_/B _7101_/B _7055_/C _7074_/A vssd1 vssd1 vccd1 vccd1 _7141_/A sky130_fd_sc_hd__a31o_1
XFILLER_101_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7065_ _7065_/A _7065_/B vssd1 vssd1 vccd1 vccd1 _7068_/A sky130_fd_sc_hd__nor2_1
XFILLER_100_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6016_ _5903_/A _6017_/B _6231_/B vssd1 vssd1 vccd1 vccd1 _6018_/A sky130_fd_sc_hd__a21o_1
XFILLER_67_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7967_ _8023_/A _7967_/B _7967_/C vssd1 vssd1 vccd1 vccd1 _8023_/B sky130_fd_sc_hd__nand3_1
X_7898_ _8207_/A _8331_/A _7898_/C _7898_/D vssd1 vssd1 vccd1 vccd1 _7948_/B sky130_fd_sc_hd__nand4_1
X_6918_ _7046_/A _7297_/B _7048_/A vssd1 vssd1 vccd1 vccd1 _6920_/B sky130_fd_sc_hd__a21oi_1
XFILLER_54_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6849_ _6942_/A _6942_/B vssd1 vssd1 vccd1 vccd1 _6970_/B sky130_fd_sc_hd__xor2_1
XFILLER_50_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8519_ _7503_/X _8716_/Q _8514_/X _8518_/X vssd1 vssd1 vccd1 vccd1 _8716_/D sky130_fd_sc_hd__o22a_1
XFILLER_2_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8749__27 vssd1 vssd1 vccd1 vccd1 _8749__27/HI _8844_/A sky130_fd_sc_hd__conb_1
XFILLER_45_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5180_ _5180_/A _5180_/B _5180_/C vssd1 vssd1 vccd1 vccd1 _5180_/X sky130_fd_sc_hd__or3_1
XFILLER_95_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8870_ _8870_/A _4387_/Y vssd1 vssd1 vccd1 vccd1 io_out[17] sky130_fd_sc_hd__ebufn_8
XFILLER_36_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7821_ _7817_/X _7651_/Y _8284_/C _7820_/Y vssd1 vssd1 vccd1 vccd1 _7822_/B sky130_fd_sc_hd__a31o_1
XFILLER_64_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7752_ _7752_/A _7752_/B _7766_/B vssd1 vssd1 vccd1 vccd1 _8111_/B sky130_fd_sc_hd__or3b_1
XFILLER_51_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4964_ _5005_/A _5007_/A _4969_/B vssd1 vssd1 vccd1 vccd1 _5076_/A sky130_fd_sc_hd__or3_1
X_8763__41 vssd1 vssd1 vccd1 vccd1 _8763__41/HI _8858_/A sky130_fd_sc_hd__conb_1
X_6703_ _6724_/A _7180_/A _6703_/C vssd1 vssd1 vccd1 vccd1 _7163_/A sky130_fd_sc_hd__nand3_1
XFILLER_32_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7683_ _7904_/A _8301_/A _7683_/C vssd1 vssd1 vccd1 vccd1 _7685_/A sky130_fd_sc_hd__and3_1
X_4895_ _5240_/A _5243_/B _5094_/A _5214_/D vssd1 vssd1 vccd1 vccd1 _4895_/X sky130_fd_sc_hd__or4_1
X_6634_ _7219_/A _7160_/B vssd1 vssd1 vccd1 vccd1 _7161_/A sky130_fd_sc_hd__nor2_1
X_6565_ _8605_/Q _8688_/Q vssd1 vssd1 vccd1 vccd1 _6566_/A sky130_fd_sc_hd__or2b_1
X_8304_ _8361_/A _8304_/B vssd1 vssd1 vccd1 vccd1 _8310_/A sky130_fd_sc_hd__xnor2_2
X_6496_ _8691_/Q vssd1 vssd1 vccd1 vccd1 _6526_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5516_ _5516_/A vssd1 vssd1 vccd1 vccd1 _5896_/A sky130_fd_sc_hd__buf_2
X_8235_ _8236_/A _8236_/B vssd1 vssd1 vccd1 vccd1 _8341_/B sky130_fd_sc_hd__or2_2
X_5447_ _5447_/A _5447_/B vssd1 vssd1 vccd1 vccd1 _5447_/X sky130_fd_sc_hd__or2_1
X_8166_ _8166_/A _8306_/A vssd1 vssd1 vccd1 vccd1 _8168_/B sky130_fd_sc_hd__or2_1
X_5378_ _8663_/Q vssd1 vssd1 vccd1 vccd1 _6371_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7117_ _7036_/A _7035_/A _7035_/B _7027_/B _7027_/A vssd1 vssd1 vccd1 vccd1 _7120_/A
+ sky130_fd_sc_hd__o32a_1
X_8097_ _8097_/A _8097_/B _8499_/A _8093_/D vssd1 vssd1 vccd1 vccd1 _8501_/A sky130_fd_sc_hd__or4bb_1
X_4329_ _4333_/A vssd1 vssd1 vccd1 vccd1 _4329_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7048_ _7048_/A _7048_/B _7048_/C vssd1 vssd1 vccd1 vccd1 _7048_/X sky130_fd_sc_hd__or3_1
XFILLER_74_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4680_ _4970_/A _4697_/B vssd1 vssd1 vccd1 vccd1 _4683_/B sky130_fd_sc_hd__nand2_1
X_6350_ _6351_/A _6364_/B vssd1 vssd1 vccd1 vccd1 _6352_/A sky130_fd_sc_hd__nor2_1
X_5301_ _8698_/Q _5285_/A _5300_/X _5296_/X vssd1 vssd1 vccd1 vccd1 _8623_/D sky130_fd_sc_hd__o211a_1
XFILLER_5_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6281_ _6186_/A _6281_/B vssd1 vssd1 vccd1 vccd1 _6281_/X sky130_fd_sc_hd__and2b_1
XFILLER_88_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8020_ _8001_/A _8020_/B vssd1 vssd1 vccd1 vccd1 _8073_/A sky130_fd_sc_hd__and2b_1
XFILLER_69_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5232_ _5105_/X _5245_/B _4937_/C _5071_/X _5092_/A vssd1 vssd1 vccd1 vccd1 _5232_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_68_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5163_ _5163_/A _5163_/B vssd1 vssd1 vccd1 vccd1 _5163_/Y sky130_fd_sc_hd__nand2_1
XFILLER_96_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5094_ _5094_/A _5094_/B vssd1 vssd1 vccd1 vccd1 _5094_/X sky130_fd_sc_hd__or2_1
X_8922_ _8922_/A _4448_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[31] sky130_fd_sc_hd__ebufn_8
X_8853_ _8853_/A _4457_/Y vssd1 vssd1 vccd1 vccd1 io_out[0] sky130_fd_sc_hd__ebufn_8
XFILLER_64_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7804_ _7804_/A _7804_/B vssd1 vssd1 vccd1 vccd1 _7805_/B sky130_fd_sc_hd__nand2_1
XFILLER_52_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5996_ _6220_/B _5996_/B vssd1 vssd1 vccd1 vccd1 _5997_/B sky130_fd_sc_hd__xnor2_1
X_7735_ _7752_/A _7747_/B vssd1 vssd1 vccd1 vccd1 _7869_/A sky130_fd_sc_hd__or2_1
X_4947_ _4985_/B vssd1 vssd1 vccd1 vccd1 _5202_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_33_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7666_ _7666_/A _7790_/A _7666_/C vssd1 vssd1 vccd1 vccd1 _7666_/X sky130_fd_sc_hd__and3_1
X_4878_ _5007_/A _5053_/D vssd1 vssd1 vccd1 vccd1 _5193_/B sky130_fd_sc_hd__or2_2
XFILLER_20_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6617_ _6617_/A _8691_/Q vssd1 vssd1 vccd1 vccd1 _6660_/A sky130_fd_sc_hd__or2b_1
XFILLER_20_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7597_ _7596_/Y _7593_/B _8535_/S vssd1 vssd1 vccd1 vccd1 _7598_/B sky130_fd_sc_hd__mux2_1
XFILLER_3_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6548_ _7540_/A _6547_/C _6628_/A vssd1 vssd1 vccd1 vccd1 _6549_/C sky130_fd_sc_hd__o21ai_1
X_6479_ _8686_/Q vssd1 vssd1 vccd1 vccd1 _7525_/A sky130_fd_sc_hd__clkbuf_1
X_8218_ _8218_/A _8327_/A _8331_/B vssd1 vssd1 vccd1 vccd1 _8218_/X sky130_fd_sc_hd__and3_1
XFILLER_87_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8149_ _8306_/A _8149_/B vssd1 vssd1 vccd1 vccd1 _8149_/Y sky130_fd_sc_hd__nand2_1
XFILLER_58_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_0 _4459_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5850_ _5850_/A _5850_/B _5850_/C vssd1 vssd1 vccd1 vccd1 _5850_/Y sky130_fd_sc_hd__nor3_1
X_4801_ _4857_/B _4898_/B vssd1 vssd1 vccd1 vccd1 _5092_/C sky130_fd_sc_hd__nor2_4
X_5781_ _5781_/A _5781_/B vssd1 vssd1 vccd1 vccd1 _5782_/B sky130_fd_sc_hd__or2_1
X_8733__11 vssd1 vssd1 vccd1 vccd1 _8733__11/HI _8828_/A sky130_fd_sc_hd__conb_1
X_7520_ _7520_/A _7520_/B vssd1 vssd1 vccd1 vccd1 _7522_/A sky130_fd_sc_hd__nor2_1
XFILLER_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4732_ _4732_/A _4732_/B _5234_/A _5224_/C vssd1 vssd1 vccd1 vccd1 _4739_/B sky130_fd_sc_hd__or4_2
X_7451_ _7395_/B _7395_/C _7395_/A vssd1 vssd1 vccd1 vccd1 _7478_/A sky130_fd_sc_hd__o21ai_1
X_4663_ _7708_/B _8594_/Q vssd1 vssd1 vccd1 vccd1 _4699_/B sky130_fd_sc_hd__and2_1
X_6402_ input2/X _8535_/S vssd1 vssd1 vccd1 vccd1 _6419_/A sky130_fd_sc_hd__and2_1
X_7382_ _7333_/A _7333_/B _7333_/C vssd1 vssd1 vccd1 vccd1 _7382_/X sky130_fd_sc_hd__o21a_1
X_4594_ _4607_/A vssd1 vssd1 vccd1 vccd1 _4639_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6333_ _6341_/A _6341_/B _6336_/A _6333_/D vssd1 vssd1 vccd1 vccd1 _6333_/X sky130_fd_sc_hd__or4_1
X_6264_ _6264_/A _6264_/B vssd1 vssd1 vccd1 vccd1 _6274_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8003_ _7948_/X _7929_/X _8020_/B _8002_/Y vssd1 vssd1 vccd1 vccd1 _8019_/A sky130_fd_sc_hd__o211ai_2
X_5215_ _5224_/C _5215_/B _5215_/C _5215_/D vssd1 vssd1 vccd1 vccd1 _5215_/X sky130_fd_sc_hd__or4_1
XFILLER_57_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6195_ _5923_/B _5973_/B _5971_/Y vssd1 vssd1 vccd1 vccd1 _6196_/A sky130_fd_sc_hd__a21oi_1
X_5146_ _4728_/A _5142_/X _5145_/X vssd1 vssd1 vccd1 vccd1 _5147_/B sky130_fd_sc_hd__o21ai_1
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5077_ _5145_/B _5256_/A vssd1 vssd1 vccd1 vccd1 _5077_/Y sky130_fd_sc_hd__nor2_1
X_8905_ _8905_/A _4428_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[14] sky130_fd_sc_hd__ebufn_8
XFILLER_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8836_ _8836_/A _4346_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[15] sky130_fd_sc_hd__ebufn_8
XFILLER_64_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5979_ _6205_/A vssd1 vssd1 vccd1 vccd1 _6269_/A sky130_fd_sc_hd__inv_2
X_7718_ _7884_/A _7862_/B vssd1 vssd1 vccd1 vccd1 _7957_/A sky130_fd_sc_hd__or2_1
XFILLER_100_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8698_ input3/X _8698_/D vssd1 vssd1 vccd1 vccd1 _8698_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7649_ _7649_/A _7654_/B vssd1 vssd1 vccd1 vccd1 _7912_/A sky130_fd_sc_hd__xnor2_2
XFILLER_4_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5000_ _5113_/A _4970_/X _4983_/X _4999_/X vssd1 vssd1 vccd1 vccd1 _5000_/X sky130_fd_sc_hd__a31o_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6951_ _6951_/A _7023_/A vssd1 vssd1 vccd1 vccd1 _6951_/X sky130_fd_sc_hd__and2_1
XFILLER_53_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6882_ _6978_/A _6866_/B _6881_/Y vssd1 vssd1 vccd1 vccd1 _6973_/A sky130_fd_sc_hd__a21oi_1
X_5902_ _5902_/A _5902_/B vssd1 vssd1 vccd1 vccd1 _5914_/A sky130_fd_sc_hd__xnor2_1
XFILLER_46_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8621_ input3/X _8621_/D vssd1 vssd1 vccd1 vccd1 _8621_/Q sky130_fd_sc_hd__dfxtp_1
X_5833_ _6044_/A _5953_/B vssd1 vssd1 vccd1 vccd1 _5954_/C sky130_fd_sc_hd__nand2_1
X_8552_ _8723_/Q _8552_/B vssd1 vssd1 vccd1 vccd1 _8556_/B sky130_fd_sc_hd__or2_1
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7503_ _7503_/A vssd1 vssd1 vccd1 vccd1 _7503_/X sky130_fd_sc_hd__clkbuf_2
X_5764_ _5764_/A _6277_/A vssd1 vssd1 vccd1 vccd1 _5764_/X sky130_fd_sc_hd__xor2_1
X_8483_ _8423_/A _8423_/B _8482_/Y vssd1 vssd1 vccd1 vccd1 _8485_/A sky130_fd_sc_hd__o21ai_1
X_5695_ _5701_/A _5695_/B vssd1 vssd1 vccd1 vccd1 _6041_/B sky130_fd_sc_hd__xnor2_1
X_4715_ _5226_/A _4716_/B vssd1 vssd1 vccd1 vccd1 _4717_/B sky130_fd_sc_hd__or2_1
X_7434_ _7434_/A _7434_/B vssd1 vssd1 vccd1 vccd1 _7446_/B sky130_fd_sc_hd__xor2_1
X_4646_ _4646_/A _4646_/B _4646_/C vssd1 vssd1 vccd1 vccd1 _4647_/A sky130_fd_sc_hd__and3_1
X_7365_ _7366_/B _7366_/C _7366_/A vssd1 vssd1 vccd1 vccd1 _7367_/A sky130_fd_sc_hd__a21oi_1
X_4577_ _8587_/Q _8590_/Q _8589_/Q vssd1 vssd1 vccd1 vccd1 _4578_/D sky130_fd_sc_hd__or3_1
X_6316_ _6316_/A _6316_/B vssd1 vssd1 vccd1 vccd1 _6316_/Y sky130_fd_sc_hd__nand2_1
XFILLER_103_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7296_ _7296_/A _7296_/B _7296_/C vssd1 vssd1 vccd1 vccd1 _7398_/A sky130_fd_sc_hd__and3_1
XFILLER_1_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6247_ _6240_/A _6240_/B _6242_/B _6242_/A _6246_/X vssd1 vssd1 vccd1 vccd1 _6298_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_57_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6178_ _6178_/A _6178_/B vssd1 vssd1 vccd1 vccd1 _6178_/X sky130_fd_sc_hd__and2_1
XFILLER_97_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5129_ _4707_/B _5001_/X _5060_/X _5128_/X vssd1 vssd1 vccd1 vccd1 _5129_/X sky130_fd_sc_hd__a31o_1
XFILLER_84_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4500_ _4810_/A vssd1 vssd1 vccd1 vccd1 _4802_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_5480_ _8600_/Q _8663_/Q vssd1 vssd1 vccd1 vccd1 _5482_/A sky130_fd_sc_hd__or2b_2
X_4431_ _4432_/A vssd1 vssd1 vccd1 vccd1 _4431_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7150_ _7151_/A _7016_/B _7149_/X vssd1 vssd1 vccd1 vccd1 _7151_/B sky130_fd_sc_hd__a21oi_1
X_4362_ _4364_/A vssd1 vssd1 vccd1 vccd1 _4362_/Y sky130_fd_sc_hd__inv_2
X_7081_ _7081_/A _7081_/B _7081_/C vssd1 vssd1 vccd1 vccd1 _7083_/A sky130_fd_sc_hd__nor3_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6101_ _6101_/A _6101_/B vssd1 vssd1 vccd1 vccd1 _6161_/B sky130_fd_sc_hd__xor2_1
XFILLER_98_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6032_ _6032_/A _6032_/B vssd1 vssd1 vccd1 vccd1 _6070_/B sky130_fd_sc_hd__xnor2_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7983_ _8021_/B _7982_/C _7982_/A vssd1 vssd1 vccd1 vccd1 _8001_/B sky130_fd_sc_hd__a21oi_1
XFILLER_66_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6934_ _6819_/A _6934_/B vssd1 vssd1 vccd1 vccd1 _6934_/X sky130_fd_sc_hd__and2b_1
XFILLER_54_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6865_ _6865_/A _7197_/B vssd1 vssd1 vccd1 vccd1 _6866_/B sky130_fd_sc_hd__xnor2_1
X_8604_ input3/X _8604_/D vssd1 vssd1 vccd1 vccd1 _8604_/Q sky130_fd_sc_hd__dfxtp_1
X_6796_ _7378_/B _7099_/A _7048_/B vssd1 vssd1 vccd1 vccd1 _6804_/A sky130_fd_sc_hd__a21oi_2
X_5816_ _5816_/A _5792_/B vssd1 vssd1 vccd1 vccd1 _5820_/A sky130_fd_sc_hd__or2b_1
X_8535_ _8534_/X _8531_/A _8535_/S vssd1 vssd1 vccd1 vccd1 _8536_/B sky130_fd_sc_hd__mux2_1
X_5747_ _5962_/A _5961_/B vssd1 vssd1 vccd1 vccd1 _5984_/A sky130_fd_sc_hd__or2b_1
XFILLER_41_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8466_ _8466_/A _8466_/B vssd1 vssd1 vccd1 vccd1 _8473_/A sky130_fd_sc_hd__xnor2_1
X_7417_ _7417_/A _7425_/B vssd1 vssd1 vccd1 vccd1 _7438_/A sky130_fd_sc_hd__xnor2_1
X_5678_ _8650_/Q _6617_/A vssd1 vssd1 vccd1 vccd1 _5679_/B sky130_fd_sc_hd__or2b_1
X_8397_ _8397_/A _8397_/B vssd1 vssd1 vccd1 vccd1 _8398_/B sky130_fd_sc_hd__xor2_1
X_4629_ _8584_/Q _8583_/Q _4623_/B _8585_/Q vssd1 vssd1 vccd1 vccd1 _4630_/C sky130_fd_sc_hd__a31o_1
X_7348_ _7348_/A _7348_/B vssd1 vssd1 vccd1 vccd1 _7390_/B sky130_fd_sc_hd__or2_1
X_7279_ _7280_/B _7279_/B vssd1 vssd1 vccd1 vccd1 _7362_/B sky130_fd_sc_hd__xnor2_1
XFILLER_103_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4980_ _5215_/B _5180_/B _5253_/C _5153_/B vssd1 vssd1 vccd1 vccd1 _4981_/D sky130_fd_sc_hd__or4_1
XFILLER_63_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6650_ _7161_/A _6651_/B vssd1 vssd1 vccd1 vccd1 _6734_/A sky130_fd_sc_hd__nand2_1
X_6581_ _6581_/A _6581_/B vssd1 vssd1 vccd1 vccd1 _6671_/A sky130_fd_sc_hd__xnor2_1
X_5601_ _5601_/A _5601_/B vssd1 vssd1 vccd1 vccd1 _5715_/B sky130_fd_sc_hd__xnor2_2
X_8320_ _8320_/A _8320_/B vssd1 vssd1 vccd1 vccd1 _8321_/B sky130_fd_sc_hd__nor2_1
X_5532_ _5513_/A _5513_/B _5531_/X vssd1 vssd1 vccd1 vccd1 _5556_/A sky130_fd_sc_hd__a21o_1
X_8251_ _8251_/A _8251_/B vssd1 vssd1 vccd1 vccd1 _8252_/B sky130_fd_sc_hd__nand2_1
X_5463_ _5463_/A _5463_/B vssd1 vssd1 vccd1 vccd1 _5475_/A sky130_fd_sc_hd__nor2_2
XFILLER_99_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7202_ _7202_/A _7258_/B vssd1 vssd1 vccd1 vccd1 _7259_/A sky130_fd_sc_hd__nand2_1
X_8182_ _8186_/A _8182_/B vssd1 vssd1 vccd1 vccd1 _8183_/B sky130_fd_sc_hd__xnor2_1
X_5394_ _8648_/Q vssd1 vssd1 vccd1 vccd1 _5414_/A sky130_fd_sc_hd__clkbuf_2
X_4414_ _4414_/A vssd1 vssd1 vccd1 vccd1 _4414_/Y sky130_fd_sc_hd__inv_2
X_7133_ _7133_/A _7133_/B vssd1 vssd1 vccd1 vccd1 _7145_/A sky130_fd_sc_hd__xnor2_2
X_4345_ _4346_/A vssd1 vssd1 vccd1 vccd1 _4345_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7064_ _7101_/C _7063_/B _7063_/C vssd1 vssd1 vccd1 vccd1 _7069_/B sky130_fd_sc_hd__a21o_1
XFILLER_74_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6015_ _6229_/A _6230_/C vssd1 vssd1 vccd1 vccd1 _6231_/B sky130_fd_sc_hd__xor2_1
XFILLER_100_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7966_ _7966_/A _7966_/B vssd1 vssd1 vccd1 vccd1 _7967_/C sky130_fd_sc_hd__xnor2_1
X_7897_ _7949_/B _7949_/C _7949_/A vssd1 vssd1 vccd1 vccd1 _7898_/D sky130_fd_sc_hd__a21o_1
X_6917_ _7048_/A _7048_/B vssd1 vssd1 vccd1 vccd1 _6920_/A sky130_fd_sc_hd__nor2_1
XFILLER_52_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6848_ _6848_/A _6848_/B vssd1 vssd1 vccd1 vccd1 _6942_/B sky130_fd_sc_hd__xnor2_2
XFILLER_50_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8518_ _8527_/A _8527_/B _8518_/C _8518_/D vssd1 vssd1 vccd1 vccd1 _8518_/X sky130_fd_sc_hd__and4_1
X_6779_ _6779_/A _6779_/B vssd1 vssd1 vccd1 vccd1 _7194_/B sky130_fd_sc_hd__xnor2_4
XFILLER_6_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8449_ _8441_/X _8442_/Y _8448_/Y vssd1 vssd1 vccd1 vccd1 _8449_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_104_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7820_ _7820_/A _7820_/B vssd1 vssd1 vccd1 vccd1 _7820_/Y sky130_fd_sc_hd__nor2_1
XFILLER_64_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7751_ _7751_/A _7751_/B vssd1 vssd1 vccd1 vccd1 _7766_/B sky130_fd_sc_hd__nor2_1
X_4963_ _5172_/B _5138_/B vssd1 vssd1 vccd1 vccd1 _4969_/B sky130_fd_sc_hd__or2_2
XFILLER_24_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6702_ _6769_/B _6702_/B vssd1 vssd1 vccd1 vccd1 _7163_/C sky130_fd_sc_hd__and2_1
X_7682_ _7682_/A _7682_/B vssd1 vssd1 vccd1 vccd1 _7683_/C sky130_fd_sc_hd__xnor2_1
X_6633_ _6645_/A vssd1 vssd1 vccd1 vccd1 _7160_/B sky130_fd_sc_hd__clkbuf_4
X_4894_ _5102_/C vssd1 vssd1 vccd1 vccd1 _5214_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_32_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6564_ _6637_/A vssd1 vssd1 vccd1 vccd1 _7425_/A sky130_fd_sc_hd__clkbuf_2
X_8303_ _8056_/B _8308_/A _8302_/X vssd1 vssd1 vccd1 vccd1 _8304_/B sky130_fd_sc_hd__o21a_1
X_6495_ _8689_/Q vssd1 vssd1 vccd1 vccd1 _6514_/A sky130_fd_sc_hd__clkbuf_2
X_5515_ _5559_/B vssd1 vssd1 vccd1 vccd1 _6082_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_8234_ _8324_/A _8324_/B vssd1 vssd1 vccd1 vccd1 _8236_/B sky130_fd_sc_hd__xnor2_1
X_5446_ _8653_/Q vssd1 vssd1 vccd1 vccd1 _5615_/A sky130_fd_sc_hd__inv_2
XFILLER_99_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8165_ _8070_/A _8070_/B _8071_/A vssd1 vssd1 vccd1 vccd1 _8178_/A sky130_fd_sc_hd__a21oi_1
X_5377_ _5376_/Y _5374_/C _7533_/B vssd1 vssd1 vccd1 vccd1 _8643_/D sky130_fd_sc_hd__a21oi_1
X_7116_ _7116_/A _7116_/B vssd1 vssd1 vccd1 vccd1 _7121_/A sky130_fd_sc_hd__xnor2_1
X_8096_ _8499_/A _8499_/B _8500_/B _8500_/A _8500_/C vssd1 vssd1 vccd1 vccd1 _8503_/B
+ sky130_fd_sc_hd__a2111o_1
X_4328_ _4459_/A vssd1 vssd1 vccd1 vccd1 _4333_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_101_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7047_ _7047_/A _7047_/B vssd1 vssd1 vccd1 vccd1 _7060_/C sky130_fd_sc_hd__xnor2_2
XFILLER_86_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7949_ _7949_/A _7949_/B _7949_/C vssd1 vssd1 vccd1 vccd1 _7949_/X sky130_fd_sc_hd__and3_1
XFILLER_70_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8809__87 vssd1 vssd1 vccd1 vccd1 _8809__87/HI _8918_/A sky130_fd_sc_hd__conb_1
XFILLER_2_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5300_ _8623_/Q _5300_/B vssd1 vssd1 vccd1 vccd1 _5300_/X sky130_fd_sc_hd__or2_1
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6280_ _6189_/A _6189_/B _6279_/X vssd1 vssd1 vccd1 vccd1 _6287_/A sky130_fd_sc_hd__a21oi_1
X_5231_ _5231_/A _5231_/B _5231_/C _5231_/D vssd1 vssd1 vccd1 vccd1 _5231_/X sky130_fd_sc_hd__or4_1
X_5162_ _5240_/A _5245_/D vssd1 vssd1 vccd1 vccd1 _5163_/B sky130_fd_sc_hd__nor2_1
XFILLER_96_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5093_ _8593_/Q _5235_/A vssd1 vssd1 vccd1 vccd1 _5166_/D sky130_fd_sc_hd__nand2_2
XFILLER_96_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8921_ _8921_/A _4447_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[30] sky130_fd_sc_hd__ebufn_8
XFILLER_49_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8852_ _8852_/A _4366_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[31] sky130_fd_sc_hd__ebufn_8
XFILLER_52_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7803_ _7804_/A _7804_/B vssd1 vssd1 vccd1 vccd1 _7936_/A sky130_fd_sc_hd__or2_1
XFILLER_37_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7734_ _8724_/Q _8600_/Q vssd1 vssd1 vccd1 vccd1 _7747_/B sky130_fd_sc_hd__and2b_1
XFILLER_52_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5995_ _5558_/A _5803_/B _5907_/B _5559_/B vssd1 vssd1 vccd1 vccd1 _5996_/B sky130_fd_sc_hd__a22oi_2
XFILLER_52_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4946_ _4946_/A _5074_/B vssd1 vssd1 vccd1 vccd1 _4985_/B sky130_fd_sc_hd__or2_1
XFILLER_33_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7665_ _7665_/A _7664_/X vssd1 vssd1 vccd1 vccd1 _7819_/A sky130_fd_sc_hd__or2b_1
X_4877_ _4959_/A _5005_/A vssd1 vssd1 vccd1 vccd1 _5053_/D sky130_fd_sc_hd__or2_2
X_6616_ _6664_/A vssd1 vssd1 vccd1 vccd1 _6657_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_7596_ _7596_/A _7596_/B vssd1 vssd1 vccd1 vccd1 _7596_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_20_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6547_ _6628_/A _7545_/B _6547_/C vssd1 vssd1 vccd1 vccd1 _6549_/B sky130_fd_sc_hd__or3_1
XFILLER_4_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6478_ _6478_/A _6478_/B _6478_/C _6478_/D vssd1 vssd1 vccd1 vccd1 _6505_/A sky130_fd_sc_hd__or4_4
X_8217_ _8406_/B vssd1 vssd1 vccd1 vccd1 _8331_/B sky130_fd_sc_hd__clkbuf_2
X_5429_ _5422_/A _5424_/Y _5428_/X vssd1 vssd1 vccd1 vccd1 _5429_/X sky130_fd_sc_hd__o21a_1
X_8148_ _8305_/B vssd1 vssd1 vccd1 vccd1 _8306_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_58_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_1 _4459_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8079_ _8079_/A _8079_/B _8079_/C vssd1 vssd1 vccd1 vccd1 _8256_/A sky130_fd_sc_hd__and3_1
XFILLER_75_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4800_ _4897_/C vssd1 vssd1 vccd1 vccd1 _4898_/B sky130_fd_sc_hd__buf_2
XFILLER_34_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5780_ _5781_/A _5781_/B vssd1 vssd1 vccd1 vccd1 _5858_/A sky130_fd_sc_hd__nand2_1
XFILLER_34_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4731_ _4731_/A vssd1 vssd1 vccd1 vccd1 _5224_/C sky130_fd_sc_hd__clkbuf_2
X_7450_ _7473_/B _7474_/B _7449_/X vssd1 vssd1 vccd1 vccd1 _7482_/B sky130_fd_sc_hd__a21oi_2
X_4662_ _4662_/A _4662_/B vssd1 vssd1 vccd1 vccd1 _4732_/B sky130_fd_sc_hd__nand2_1
X_6401_ _6406_/B _7552_/A vssd1 vssd1 vccd1 vccd1 _8535_/S sky130_fd_sc_hd__or2_4
X_7381_ _7397_/A _7397_/B vssd1 vssd1 vccd1 vccd1 _7381_/Y sky130_fd_sc_hd__nand2_1
X_4593_ _8574_/Q _4598_/C vssd1 vssd1 vccd1 vccd1 _4597_/A sky130_fd_sc_hd__and2_1
X_6332_ _6332_/A _6332_/B vssd1 vssd1 vccd1 vccd1 _6333_/D sky130_fd_sc_hd__nor2_1
X_6263_ _6263_/A _6263_/B vssd1 vssd1 vccd1 vccd1 _6264_/B sky130_fd_sc_hd__xnor2_2
X_8002_ _8001_/A _8001_/B _8001_/C vssd1 vssd1 vccd1 vccd1 _8002_/Y sky130_fd_sc_hd__o21ai_1
X_5214_ _5214_/A _5214_/B _5214_/C _5214_/D vssd1 vssd1 vccd1 vccd1 _5214_/X sky130_fd_sc_hd__or4_1
X_6194_ _6292_/B _6194_/B vssd1 vssd1 vccd1 vccd1 _6197_/A sky130_fd_sc_hd__xnor2_2
XFILLER_84_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5145_ _5190_/B _5145_/B _5149_/B _5149_/D vssd1 vssd1 vccd1 vccd1 _5145_/X sky130_fd_sc_hd__or4_1
XFILLER_84_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5076_ _5076_/A vssd1 vssd1 vccd1 vccd1 _5256_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_8904_ _8904_/A _4425_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[13] sky130_fd_sc_hd__ebufn_8
XFILLER_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8835_ _8835_/A _4345_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[14] sky130_fd_sc_hd__ebufn_8
XFILLER_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5978_ _5918_/A _5918_/B _5977_/X vssd1 vssd1 vccd1 vccd1 _6024_/A sky130_fd_sc_hd__a21oi_1
X_8697_ input3/X _8697_/D vssd1 vssd1 vccd1 vccd1 _8697_/Q sky130_fd_sc_hd__dfxtp_1
X_7717_ _7717_/A _7717_/B vssd1 vssd1 vccd1 vccd1 _7862_/B sky130_fd_sc_hd__xnor2_2
XFILLER_12_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4929_ _5083_/A vssd1 vssd1 vccd1 vccd1 _4990_/A sky130_fd_sc_hd__clkbuf_2
X_7648_ _8051_/A vssd1 vssd1 vccd1 vccd1 _7666_/A sky130_fd_sc_hd__clkbuf_2
X_7579_ _8708_/Q vssd1 vssd1 vccd1 vccd1 _7627_/A sky130_fd_sc_hd__clkinv_2
XFILLER_85_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6950_ _6950_/A _6950_/B vssd1 vssd1 vccd1 vccd1 _7039_/A sky130_fd_sc_hd__xnor2_2
XFILLER_66_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5901_ _5901_/A _5900_/X vssd1 vssd1 vccd1 vccd1 _5902_/B sky130_fd_sc_hd__or2b_1
X_6881_ _6881_/A _7197_/B vssd1 vssd1 vccd1 vccd1 _6881_/Y sky130_fd_sc_hd__nor2_1
X_8620_ input3/X _8620_/D vssd1 vssd1 vccd1 vccd1 _8620_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5832_ _5832_/A vssd1 vssd1 vccd1 vccd1 _5954_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_34_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8551_ _8566_/A _8552_/B vssd1 vssd1 vccd1 vccd1 _8556_/A sky130_fd_sc_hd__nand2_1
X_5763_ _5763_/A _5828_/A vssd1 vssd1 vccd1 vccd1 _6277_/A sky130_fd_sc_hd__xnor2_4
XFILLER_22_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7502_ _6334_/X _8696_/Q _7498_/Y _7501_/Y vssd1 vssd1 vccd1 vccd1 _8696_/D sky130_fd_sc_hd__o22a_1
X_4714_ _6777_/B vssd1 vssd1 vccd1 vccd1 _5226_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_8482_ _8482_/A _8482_/B vssd1 vssd1 vccd1 vccd1 _8482_/Y sky130_fd_sc_hd__nand2_1
X_5694_ _6046_/A _6046_/B _5693_/X vssd1 vssd1 vccd1 vccd1 _6051_/B sky130_fd_sc_hd__a21oi_2
XFILLER_30_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7433_ _7433_/A vssd1 vssd1 vccd1 vccd1 _7436_/B sky130_fd_sc_hd__inv_2
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4645_ _8590_/Q _4645_/B vssd1 vssd1 vccd1 vccd1 _4646_/C sky130_fd_sc_hd__nand2_2
X_7364_ _7456_/A _7455_/B vssd1 vssd1 vccd1 vccd1 _7366_/A sky130_fd_sc_hd__xnor2_1
X_4576_ _8586_/Q _8585_/Q _8588_/Q _8591_/Q vssd1 vssd1 vccd1 vccd1 _4578_/C sky130_fd_sc_hd__or4b_1
X_6315_ _6316_/A _6316_/B vssd1 vssd1 vccd1 vccd1 _6315_/X sky130_fd_sc_hd__or2_1
X_7295_ _7439_/A _7378_/B _7378_/D vssd1 vssd1 vccd1 vccd1 _7327_/A sky130_fd_sc_hd__or3b_1
X_6246_ _6241_/A _6246_/B vssd1 vssd1 vccd1 vccd1 _6246_/X sky130_fd_sc_hd__and2b_1
XFILLER_39_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6177_ _5990_/A _5990_/B _5991_/B _5991_/A vssd1 vssd1 vccd1 vccd1 _6292_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_57_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5128_ _4953_/X _5190_/A _5082_/X _5126_/X _5261_/A vssd1 vssd1 vccd1 vccd1 _5128_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5059_ _5066_/A _5050_/Y _5058_/Y _4953_/A vssd1 vssd1 vccd1 vccd1 _5059_/X sky130_fd_sc_hd__a211o_1
XFILLER_44_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4430_ _4432_/A vssd1 vssd1 vccd1 vccd1 _4430_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4361_ _4364_/A vssd1 vssd1 vccd1 vccd1 _4361_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6100_ _6157_/A _6157_/B _6099_/Y vssd1 vssd1 vccd1 vccd1 _6161_/A sky130_fd_sc_hd__o21a_1
X_7080_ _6964_/B _6964_/C _6964_/A vssd1 vssd1 vccd1 vccd1 _7081_/C sky130_fd_sc_hd__o21ba_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6031_ _6317_/A _6244_/B vssd1 vssd1 vccd1 vccd1 _6306_/A sky130_fd_sc_hd__and2_1
XFILLER_100_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7982_ _7982_/A _8021_/B _7982_/C vssd1 vssd1 vccd1 vccd1 _8001_/A sky130_fd_sc_hd__and3_1
XFILLER_66_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6933_ _6932_/A _6932_/B _6932_/C vssd1 vssd1 vccd1 vccd1 _6936_/B sky130_fd_sc_hd__a21o_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6864_ _6864_/A vssd1 vssd1 vccd1 vccd1 _7197_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_62_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8603_ input3/X _8603_/D vssd1 vssd1 vccd1 vccd1 _8603_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5815_ _5815_/A _5877_/B vssd1 vssd1 vccd1 vccd1 _5822_/A sky130_fd_sc_hd__xnor2_2
X_6795_ _7067_/A vssd1 vssd1 vccd1 vccd1 _7099_/A sky130_fd_sc_hd__clkbuf_2
X_8534_ _8532_/Y _8534_/B vssd1 vssd1 vccd1 vccd1 _8534_/X sky130_fd_sc_hd__and2b_1
X_5746_ _5746_/A _5746_/B vssd1 vssd1 vccd1 vccd1 _5768_/A sky130_fd_sc_hd__nand2_1
XFILLER_22_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8465_ _8465_/A _8465_/B vssd1 vssd1 vccd1 vccd1 _8466_/B sky130_fd_sc_hd__xnor2_1
X_5677_ _6042_/B vssd1 vssd1 vccd1 vccd1 _6180_/A sky130_fd_sc_hd__clkbuf_2
X_7416_ _7416_/A _7416_/B vssd1 vssd1 vccd1 vccd1 _7428_/A sky130_fd_sc_hd__xor2_1
X_4628_ _8584_/Q _8585_/Q _4628_/C vssd1 vssd1 vccd1 vccd1 _4632_/B sky130_fd_sc_hd__and3_1
X_8396_ _8462_/A _8396_/B vssd1 vssd1 vccd1 vccd1 _8397_/B sky130_fd_sc_hd__nor2_1
XFILLER_104_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7347_ _7345_/X _7344_/Y _7333_/Y _7333_/A vssd1 vssd1 vccd1 vccd1 _7348_/B sky130_fd_sc_hd__a211oi_1
X_4559_ _8623_/Q _4563_/B vssd1 vssd1 vccd1 vccd1 _4560_/A sky130_fd_sc_hd__and2_1
XFILLER_1_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7278_ _7278_/A _7278_/B vssd1 vssd1 vccd1 vccd1 _7279_/B sky130_fd_sc_hd__xnor2_1
XFILLER_89_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6229_ _6229_/A vssd1 vssd1 vccd1 vccd1 _6230_/B sky130_fd_sc_hd__clkinv_2
XFILLER_57_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8784__62 vssd1 vssd1 vccd1 vccd1 _8784__62/HI _8893_/A sky130_fd_sc_hd__conb_1
XFILLER_82_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6580_ _6591_/A _6580_/B vssd1 vssd1 vccd1 vccd1 _7175_/A sky130_fd_sc_hd__xnor2_2
X_5600_ _5600_/A _5600_/B vssd1 vssd1 vccd1 vccd1 _5601_/B sky130_fd_sc_hd__xnor2_2
X_5531_ _6214_/A _5531_/B vssd1 vssd1 vccd1 vccd1 _5531_/X sky130_fd_sc_hd__and2_1
X_8250_ _8251_/A _8251_/B vssd1 vssd1 vccd1 vccd1 _8298_/A sky130_fd_sc_hd__nor2_1
X_7201_ _6876_/C _7192_/Y _7200_/Y vssd1 vssd1 vccd1 vccd1 _7258_/B sky130_fd_sc_hd__a21bo_1
X_5462_ _8597_/Q _5462_/B vssd1 vssd1 vccd1 vccd1 _5463_/B sky130_fd_sc_hd__and2b_1
X_8181_ _8181_/A _8181_/B vssd1 vssd1 vccd1 vccd1 _8182_/B sky130_fd_sc_hd__xor2_1
X_4413_ _4414_/A vssd1 vssd1 vccd1 vccd1 _4413_/Y sky130_fd_sc_hd__inv_2
X_5393_ _8651_/Q vssd1 vssd1 vccd1 vccd1 _5447_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7132_ _7132_/A _7132_/B vssd1 vssd1 vccd1 vccd1 _7133_/B sky130_fd_sc_hd__xnor2_1
X_4344_ _4346_/A vssd1 vssd1 vccd1 vccd1 _4344_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7063_ _7101_/C _7063_/B _7063_/C vssd1 vssd1 vccd1 vccd1 _7101_/D sky130_fd_sc_hd__nand3_2
XFILLER_98_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6014_ _6224_/A _6014_/B vssd1 vssd1 vccd1 vccd1 _6230_/C sky130_fd_sc_hd__xnor2_1
XFILLER_100_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7965_ _8395_/A _8134_/B _7964_/X vssd1 vssd1 vccd1 vccd1 _7966_/B sky130_fd_sc_hd__a21oi_1
XFILLER_82_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7896_ _7949_/A _7949_/B _7949_/C vssd1 vssd1 vccd1 vccd1 _7898_/C sky130_fd_sc_hd__nand3_1
X_6916_ _7418_/A _7239_/A vssd1 vssd1 vccd1 vccd1 _6922_/A sky130_fd_sc_hd__nor2_1
XFILLER_35_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6847_ _6847_/A _7092_/C vssd1 vssd1 vccd1 vccd1 _6848_/B sky130_fd_sc_hd__xor2_2
XFILLER_22_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6778_ _6778_/A _6778_/B vssd1 vssd1 vccd1 vccd1 _6779_/B sky130_fd_sc_hd__nor2_2
XFILLER_52_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8517_ _8520_/A _8520_/B vssd1 vssd1 vccd1 vccd1 _8518_/D sky130_fd_sc_hd__nand2_1
X_5729_ _5742_/A _5729_/B vssd1 vssd1 vccd1 vccd1 _5789_/B sky130_fd_sc_hd__xnor2_1
XFILLER_50_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8448_ _8448_/A _8448_/B vssd1 vssd1 vccd1 vccd1 _8448_/Y sky130_fd_sc_hd__xnor2_1
X_8379_ _8385_/A _8379_/B vssd1 vssd1 vccd1 vccd1 _8390_/A sky130_fd_sc_hd__nor2_1
XFILLER_104_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7750_ _7871_/A _8725_/Q vssd1 vssd1 vccd1 vccd1 _7751_/B sky130_fd_sc_hd__and2b_1
X_4962_ _5054_/C _5180_/B vssd1 vssd1 vccd1 vccd1 _5138_/B sky130_fd_sc_hd__or2_2
X_6701_ _6700_/B _6673_/A _6685_/A vssd1 vssd1 vccd1 vccd1 _6702_/B sky130_fd_sc_hd__a21o_1
X_7681_ _7912_/A _8305_/A vssd1 vssd1 vccd1 vccd1 _7682_/B sky130_fd_sc_hd__nor2_1
X_4893_ _5046_/A _5122_/A vssd1 vssd1 vccd1 vccd1 _5102_/C sky130_fd_sc_hd__or2_2
XFILLER_32_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6632_ _7296_/A _6639_/A _6794_/A vssd1 vssd1 vccd1 vccd1 _6645_/A sky130_fd_sc_hd__mux2_1
X_6563_ _6844_/A vssd1 vssd1 vccd1 vccd1 _6637_/A sky130_fd_sc_hd__inv_2
X_8302_ _8302_/A _8446_/S vssd1 vssd1 vccd1 vccd1 _8302_/X sky130_fd_sc_hd__or2_1
X_5514_ _5514_/A _5526_/C vssd1 vssd1 vccd1 vccd1 _6033_/A sky130_fd_sc_hd__xnor2_1
X_6494_ _8690_/Q vssd1 vssd1 vccd1 vccd1 _6520_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_8233_ _8337_/B _8233_/B vssd1 vssd1 vccd1 vccd1 _8324_/B sky130_fd_sc_hd__nand2_1
X_5445_ _5413_/X _5444_/X _5441_/A _4582_/B vssd1 vssd1 vccd1 vccd1 _8652_/D sky130_fd_sc_hd__o2bb2a_1
X_8164_ _8189_/A _8164_/B vssd1 vssd1 vccd1 vccd1 _8181_/A sky130_fd_sc_hd__xnor2_1
X_7115_ _7051_/B _7115_/B vssd1 vssd1 vccd1 vccd1 _7116_/B sky130_fd_sc_hd__and2b_1
X_5376_ _8643_/Q vssd1 vssd1 vccd1 vccd1 _5376_/Y sky130_fd_sc_hd__inv_2
X_4327_ _4451_/A vssd1 vssd1 vccd1 vccd1 _4459_/A sky130_fd_sc_hd__buf_6
X_8095_ _8499_/A _8093_/D _8097_/A _8097_/B vssd1 vssd1 vccd1 vccd1 _8500_/C sky130_fd_sc_hd__o2bb2a_1
XFILLER_59_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7046_ _7046_/A _7245_/B vssd1 vssd1 vccd1 vccd1 _7047_/B sky130_fd_sc_hd__xnor2_1
XFILLER_101_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7948_ _7948_/A _7948_/B _7948_/C vssd1 vssd1 vccd1 vccd1 _7948_/X sky130_fd_sc_hd__and3_1
XFILLER_70_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8754__32 vssd1 vssd1 vccd1 vccd1 _8754__32/HI _8849_/A sky130_fd_sc_hd__conb_1
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7879_ _7879_/A _7879_/B vssd1 vssd1 vccd1 vccd1 _7880_/C sky130_fd_sc_hd__xor2_2
XFILLER_10_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5230_ _5230_/A _5230_/B _5230_/C vssd1 vssd1 vccd1 vccd1 _5230_/X sky130_fd_sc_hd__and3_1
XFILLER_69_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5161_ _5138_/B _5199_/A _5149_/X _5160_/X _5060_/A vssd1 vssd1 vccd1 vccd1 _5161_/X
+ sky130_fd_sc_hd__o311a_1
X_5092_ _5092_/A _5231_/C _5092_/C _5231_/D vssd1 vssd1 vccd1 vccd1 _5215_/D sky130_fd_sc_hd__or4_1
X_8920_ _8920_/A _4446_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[29] sky130_fd_sc_hd__ebufn_8
XFILLER_83_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8851_ _8851_/A _4364_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[30] sky130_fd_sc_hd__ebufn_8
X_7802_ _7664_/X _7685_/X _7924_/B vssd1 vssd1 vccd1 vccd1 _7804_/B sky130_fd_sc_hd__a21bo_1
XFILLER_64_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5994_ _5902_/A _5900_/X _5901_/A vssd1 vssd1 vccd1 vccd1 _5998_/A sky130_fd_sc_hd__a21o_1
X_7733_ _6608_/B _8724_/Q vssd1 vssd1 vccd1 vccd1 _7752_/A sky130_fd_sc_hd__and2b_1
X_4945_ _5122_/A _4969_/C vssd1 vssd1 vccd1 vccd1 _5176_/B sky130_fd_sc_hd__or2_1
XFILLER_24_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7664_ _7664_/A _7790_/A _7995_/B _8050_/A vssd1 vssd1 vccd1 vccd1 _7664_/X sky130_fd_sc_hd__or4b_1
X_4876_ _5041_/B _4898_/B vssd1 vssd1 vccd1 vccd1 _5005_/A sky130_fd_sc_hd__nor2_1
XFILLER_20_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7595_ _7627_/A _7589_/B _7588_/A vssd1 vssd1 vccd1 vccd1 _7596_/B sky130_fd_sc_hd__o21a_1
X_6615_ _7676_/A _6539_/A vssd1 vssd1 vccd1 vccd1 _6664_/A sky130_fd_sc_hd__or2b_1
X_6546_ _6536_/A _6533_/C _6540_/D _6545_/X vssd1 vssd1 vccd1 vccd1 _6547_/C sky130_fd_sc_hd__o31a_1
X_6477_ _6477_/A _6477_/B _6477_/C vssd1 vssd1 vccd1 vccd1 _6478_/D sky130_fd_sc_hd__or3_1
X_8216_ _7752_/A _7751_/B _7752_/B _7875_/X _7746_/A vssd1 vssd1 vccd1 vccd1 _8406_/B
+ sky130_fd_sc_hd__o311a_1
X_5428_ _5428_/A _8646_/Q vssd1 vssd1 vccd1 vccd1 _5428_/X sky130_fd_sc_hd__xor2_1
XFILLER_99_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8147_ _8147_/A _8302_/A vssd1 vssd1 vccd1 vccd1 _8149_/B sky130_fd_sc_hd__nor2_1
X_5359_ _5359_/A _5359_/B vssd1 vssd1 vccd1 vccd1 _8637_/D sky130_fd_sc_hd__nor2_1
X_8078_ _8057_/A _7996_/A _8147_/A vssd1 vssd1 vccd1 vccd1 _8079_/C sky130_fd_sc_hd__o21a_1
XFILLER_58_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_2 _4459_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7029_ _7092_/C _7114_/B vssd1 vssd1 vccd1 vccd1 _7034_/A sky130_fd_sc_hd__xnor2_1
XFILLER_82_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4730_ _5135_/A _4989_/A vssd1 vssd1 vccd1 vccd1 _4731_/A sky130_fd_sc_hd__nand2_1
X_4661_ _4661_/A _4739_/A vssd1 vssd1 vccd1 vccd1 _4697_/B sky130_fd_sc_hd__nand2_1
X_7380_ _7380_/A _7380_/B vssd1 vssd1 vccd1 vccd1 _7397_/B sky130_fd_sc_hd__xnor2_1
X_6400_ _6400_/A _6400_/B _6400_/C vssd1 vssd1 vccd1 vccd1 _7552_/A sky130_fd_sc_hd__and3_2
X_4592_ _4592_/A vssd1 vssd1 vccd1 vccd1 _8573_/D sky130_fd_sc_hd__clkbuf_1
X_6331_ _6332_/A _6332_/B vssd1 vssd1 vccd1 vccd1 _6336_/A sky130_fd_sc_hd__and2_1
XFILLER_6_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6262_ _6262_/A _6262_/B vssd1 vssd1 vccd1 vccd1 _6263_/B sky130_fd_sc_hd__xnor2_1
X_8001_ _8001_/A _8001_/B _8001_/C vssd1 vssd1 vccd1 vccd1 _8020_/B sky130_fd_sc_hd__or3_1
X_6193_ _6193_/A _6193_/B vssd1 vssd1 vccd1 vccd1 _6194_/B sky130_fd_sc_hd__xnor2_1
X_5213_ _5213_/A _5213_/B _5213_/C vssd1 vssd1 vccd1 vccd1 _5213_/X sky130_fd_sc_hd__and3_1
X_5144_ _5159_/A _5144_/B vssd1 vssd1 vccd1 vccd1 _5149_/D sky130_fd_sc_hd__nand2_1
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5075_ _5143_/A _5075_/B vssd1 vssd1 vccd1 vccd1 _5075_/Y sky130_fd_sc_hd__nor2_1
X_8903_ _8903_/A _4423_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[12] sky130_fd_sc_hd__ebufn_8
X_8834_ _8834_/A _4344_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[13] sky130_fd_sc_hd__ebufn_8
XFILLER_25_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5977_ _5917_/A _5977_/B vssd1 vssd1 vccd1 vccd1 _5977_/X sky130_fd_sc_hd__and2b_1
X_8696_ input3/X _8696_/D vssd1 vssd1 vccd1 vccd1 _8696_/Q sky130_fd_sc_hd__dfxtp_1
X_7716_ _7745_/A _7745_/B _7693_/A vssd1 vssd1 vccd1 vccd1 _7717_/A sky130_fd_sc_hd__a21o_1
X_4928_ _4928_/A _4928_/B vssd1 vssd1 vccd1 vccd1 _4928_/Y sky130_fd_sc_hd__nand2_1
XFILLER_40_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7647_ _7986_/A vssd1 vssd1 vccd1 vccd1 _8051_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4859_ _4859_/A _4898_/A vssd1 vssd1 vccd1 vccd1 _5119_/B sky130_fd_sc_hd__nor2_1
X_7578_ _7615_/B _7552_/Y _7575_/Y _7577_/X _7541_/X vssd1 vssd1 vccd1 vccd1 _8707_/D
+ sky130_fd_sc_hd__a221o_1
X_6529_ _6529_/A _6529_/B vssd1 vssd1 vccd1 vccd1 _6529_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_79_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5900_ _5900_/A _5900_/B _5900_/C vssd1 vssd1 vccd1 vccd1 _5900_/X sky130_fd_sc_hd__or3_1
X_6880_ _6880_/A _6880_/B vssd1 vssd1 vccd1 vccd1 _6887_/A sky130_fd_sc_hd__and2_1
XFILLER_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5831_ _5831_/A _5831_/B vssd1 vssd1 vccd1 vccd1 _5838_/A sky130_fd_sc_hd__xor2_1
X_8550_ _8546_/A _6427_/X _8549_/X vssd1 vssd1 vccd1 vccd1 _8722_/D sky130_fd_sc_hd__a21bo_1
X_5762_ _6185_/A vssd1 vssd1 vccd1 vccd1 _5828_/A sky130_fd_sc_hd__clkinv_2
X_7501_ _7509_/A _7501_/B vssd1 vssd1 vccd1 vccd1 _7501_/Y sky130_fd_sc_hd__nor2_1
X_4713_ _4713_/A vssd1 vssd1 vccd1 vccd1 _8598_/D sky130_fd_sc_hd__clkbuf_1
X_8481_ _8481_/A _8481_/B vssd1 vssd1 vccd1 vccd1 _8486_/A sky130_fd_sc_hd__xnor2_1
X_5693_ _5922_/A _5701_/A _5749_/B vssd1 vssd1 vccd1 vccd1 _5693_/X sky130_fd_sc_hd__and3_1
XFILLER_30_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7432_ _7417_/A _7231_/A _7403_/X vssd1 vssd1 vccd1 vccd1 _7433_/A sky130_fd_sc_hd__a21o_1
X_4644_ _8590_/Q _4645_/B vssd1 vssd1 vccd1 vccd1 _4646_/B sky130_fd_sc_hd__or2_1
X_7363_ _7454_/A _7363_/B vssd1 vssd1 vccd1 vccd1 _7455_/B sky130_fd_sc_hd__xnor2_1
X_4575_ _8574_/Q _8573_/Q _8576_/Q _8575_/Q vssd1 vssd1 vccd1 vccd1 _4578_/B sky130_fd_sc_hd__or4_1
XFILLER_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7294_ _7294_/A _7294_/B vssd1 vssd1 vccd1 vccd1 _7378_/D sky130_fd_sc_hd__xnor2_1
X_6314_ _6314_/A _6314_/B vssd1 vssd1 vccd1 vccd1 _6314_/Y sky130_fd_sc_hd__nor2_1
X_6245_ _6306_/A _6306_/B _6317_/B _6244_/Y _6243_/B vssd1 vssd1 vccd1 vccd1 _6299_/A
+ sky130_fd_sc_hd__a32o_2
X_6176_ _6025_/A _6025_/B _6175_/X vssd1 vssd1 vccd1 vccd1 _6240_/A sky130_fd_sc_hd__a21o_1
X_5127_ _5127_/A _5127_/B vssd1 vssd1 vccd1 vccd1 _5261_/A sky130_fd_sc_hd__or2_1
X_5058_ _5173_/B _5058_/B vssd1 vssd1 vccd1 vccd1 _5058_/Y sky130_fd_sc_hd__nor2_1
XFILLER_72_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8679_ input3/X _8679_/D vssd1 vssd1 vccd1 vccd1 _8679_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4360_ _4364_/A vssd1 vssd1 vccd1 vccd1 _4360_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6030_ _6075_/A _6030_/B vssd1 vssd1 vccd1 vccd1 _6244_/B sky130_fd_sc_hd__nand2_1
XFILLER_66_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7981_ _8021_/A _7980_/C _7980_/A vssd1 vssd1 vccd1 vccd1 _7982_/C sky130_fd_sc_hd__a21o_1
XFILLER_66_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6932_ _6932_/A _6932_/B _6932_/C vssd1 vssd1 vccd1 vccd1 _6936_/A sky130_fd_sc_hd__nand3_1
XFILLER_54_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6863_ _6863_/A _6869_/A vssd1 vssd1 vccd1 vccd1 _6865_/A sky130_fd_sc_hd__nor2_1
XFILLER_81_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8602_ input3/X _8602_/D vssd1 vssd1 vccd1 vccd1 _8602_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5814_ _5814_/A _5814_/B vssd1 vssd1 vccd1 vccd1 _5877_/B sky130_fd_sc_hd__xnor2_2
X_6794_ _6794_/A _6814_/A vssd1 vssd1 vccd1 vccd1 _7067_/A sky130_fd_sc_hd__xnor2_1
XFILLER_10_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8533_ _8533_/A _8533_/B vssd1 vssd1 vccd1 vccd1 _8534_/B sky130_fd_sc_hd__nand2_1
X_5745_ _5745_/A _5786_/B vssd1 vssd1 vccd1 vccd1 _5770_/A sky130_fd_sc_hd__xnor2_1
X_8464_ _8464_/A _8464_/B vssd1 vssd1 vccd1 vccd1 _8465_/B sky130_fd_sc_hd__xnor2_1
X_5676_ _5746_/A _5746_/B vssd1 vssd1 vccd1 vccd1 _5688_/A sky130_fd_sc_hd__xnor2_1
X_7415_ _7413_/A _7412_/C _7412_/B vssd1 vssd1 vccd1 vccd1 _7449_/B sky130_fd_sc_hd__a21o_1
X_4627_ _8584_/Q _4628_/C _4626_/Y vssd1 vssd1 vccd1 vccd1 _8584_/D sky130_fd_sc_hd__a21oi_1
X_8395_ _8395_/A _8395_/B vssd1 vssd1 vccd1 vccd1 _8396_/B sky130_fd_sc_hd__xnor2_1
X_4558_ _4558_/A vssd1 vssd1 vccd1 vccd1 _8876_/A sky130_fd_sc_hd__clkbuf_1
X_7346_ _7333_/A _7333_/Y _7344_/Y _7345_/X vssd1 vssd1 vccd1 vccd1 _7348_/A sky130_fd_sc_hd__o211a_1
XFILLER_89_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7277_ _7353_/A _7353_/B _7276_/Y vssd1 vssd1 vccd1 vccd1 _7280_/B sky130_fd_sc_hd__a21o_1
XFILLER_89_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4489_ _6617_/A vssd1 vssd1 vccd1 vccd1 _4820_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6228_ _6228_/A _6228_/B vssd1 vssd1 vccd1 vccd1 _6233_/A sky130_fd_sc_hd__xor2_2
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6159_ _6304_/B _6159_/B vssd1 vssd1 vccd1 vccd1 _6316_/B sky130_fd_sc_hd__xnor2_1
XFILLER_85_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5530_ _5993_/A _6009_/A vssd1 vssd1 vccd1 vccd1 _6214_/A sky130_fd_sc_hd__nor2_4
X_5461_ _5462_/B _8597_/Q vssd1 vssd1 vccd1 vccd1 _5463_/A sky130_fd_sc_hd__and2b_1
X_7200_ _7234_/A _7234_/B vssd1 vssd1 vccd1 vccd1 _7200_/Y sky130_fd_sc_hd__nand2_1
X_4412_ _4414_/A vssd1 vssd1 vccd1 vccd1 _4412_/Y sky130_fd_sc_hd__inv_2
X_8180_ _8180_/A _8180_/B vssd1 vssd1 vccd1 vccd1 _8181_/B sky130_fd_sc_hd__xor2_1
X_5392_ _8652_/Q vssd1 vssd1 vccd1 vccd1 _5441_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7131_ _7131_/A _7131_/B vssd1 vssd1 vccd1 vccd1 _7132_/B sky130_fd_sc_hd__xnor2_1
X_4343_ _4346_/A vssd1 vssd1 vccd1 vccd1 _4343_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7062_ _7062_/A _7062_/B vssd1 vssd1 vccd1 vccd1 _7063_/C sky130_fd_sc_hd__nand2_1
XFILLER_86_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6013_ _6013_/A _6013_/B vssd1 vssd1 vccd1 vccd1 _6019_/A sky130_fd_sc_hd__nor2_1
XFILLER_94_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7964_ _7964_/A vssd1 vssd1 vccd1 vccd1 _7964_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_82_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6915_ _6914_/A _6914_/B _6914_/C vssd1 vssd1 vccd1 vccd1 _7044_/B sky130_fd_sc_hd__a21oi_1
X_7895_ _7894_/A _7894_/B _7894_/C vssd1 vssd1 vccd1 vccd1 _7949_/C sky130_fd_sc_hd__a21o_1
X_6846_ _6751_/A _6831_/B _7088_/A vssd1 vssd1 vccd1 vccd1 _7092_/C sky130_fd_sc_hd__a21bo_2
X_6777_ _7533_/A _6777_/B vssd1 vssd1 vccd1 vccd1 _6778_/A sky130_fd_sc_hd__nor2_1
X_8516_ _8520_/A _8520_/B vssd1 vssd1 vccd1 vccd1 _8518_/C sky130_fd_sc_hd__or2_1
X_5728_ _5792_/A _5792_/B vssd1 vssd1 vccd1 vccd1 _5729_/B sky130_fd_sc_hd__xor2_1
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8447_ _8447_/A _8447_/B vssd1 vssd1 vccd1 vccd1 _8448_/B sky130_fd_sc_hd__xnor2_1
X_5659_ _5826_/A _5922_/A vssd1 vssd1 vccd1 vccd1 _5659_/Y sky130_fd_sc_hd__nand2_1
X_8378_ _8376_/Y _8345_/B _8377_/Y vssd1 vssd1 vccd1 vccd1 _8435_/A sky130_fd_sc_hd__a21o_1
XFILLER_104_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7329_ _7325_/B _7325_/C _7325_/A vssd1 vssd1 vccd1 vccd1 _7330_/C sky130_fd_sc_hd__a21o_1
XFILLER_77_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4961_ _4961_/A _4961_/B vssd1 vssd1 vccd1 vccd1 _5180_/B sky130_fd_sc_hd__nor2_2
X_6700_ _6719_/A _6700_/B _6769_/A vssd1 vssd1 vccd1 vccd1 _6769_/B sky130_fd_sc_hd__nand3_1
X_7680_ _7789_/A _7789_/B vssd1 vssd1 vccd1 vccd1 _8301_/A sky130_fd_sc_hd__xnor2_4
X_4892_ _5026_/A _5227_/B _5026_/B vssd1 vssd1 vccd1 vccd1 _5122_/A sky130_fd_sc_hd__and3_1
X_6631_ _6614_/X _6657_/B _6657_/C _6629_/A _7175_/A vssd1 vssd1 vccd1 vccd1 _6794_/A
+ sky130_fd_sc_hd__a311o_1
X_8301_ _8301_/A _8301_/B vssd1 vssd1 vccd1 vccd1 _8308_/A sky130_fd_sc_hd__and2_1
X_6562_ _6562_/A _6562_/B vssd1 vssd1 vccd1 vccd1 _6844_/A sky130_fd_sc_hd__xnor2_4
X_5513_ _5513_/A _5513_/B vssd1 vssd1 vccd1 vccd1 _5526_/C sky130_fd_sc_hd__xor2_1
X_6493_ _8692_/Q vssd1 vssd1 vccd1 vccd1 _6536_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_8232_ _8232_/A _8410_/B vssd1 vssd1 vccd1 vccd1 _8233_/B sky130_fd_sc_hd__nand2_1
X_5444_ _5444_/A _5444_/B vssd1 vssd1 vccd1 vccd1 _5444_/X sky130_fd_sc_hd__or2_1
XFILLER_99_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8163_ _8163_/A _8163_/B vssd1 vssd1 vccd1 vccd1 _8164_/B sky130_fd_sc_hd__xor2_1
X_7114_ _7265_/A _7114_/B vssd1 vssd1 vccd1 vccd1 _7116_/A sky130_fd_sc_hd__nor2_1
X_5375_ _5375_/A vssd1 vssd1 vccd1 vccd1 _8642_/D sky130_fd_sc_hd__clkbuf_1
X_4326_ input1/X vssd1 vssd1 vccd1 vccd1 _4451_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_8094_ _8094_/A _8097_/B vssd1 vssd1 vccd1 vccd1 _8500_/A sky130_fd_sc_hd__or2_1
XFILLER_59_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7045_ _7045_/A _7045_/B vssd1 vssd1 vccd1 vccd1 _7051_/B sky130_fd_sc_hd__nor2_1
XFILLER_101_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7947_ _7847_/Y _8522_/A _7946_/X vssd1 vssd1 vccd1 vccd1 _8527_/A sky130_fd_sc_hd__a21o_1
XFILLER_27_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7878_ _8218_/A _7964_/A _7877_/Y vssd1 vssd1 vccd1 vccd1 _7879_/B sky130_fd_sc_hd__a21oi_2
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6829_ _6766_/A _6829_/B vssd1 vssd1 vccd1 vccd1 _6829_/X sky130_fd_sc_hd__and2b_1
XFILLER_23_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5160_ _5155_/X _5159_/X _4953_/X vssd1 vssd1 vccd1 vccd1 _5160_/X sky130_fd_sc_hd__a21o_1
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5091_ _5091_/A _5098_/B _5215_/C _5091_/D vssd1 vssd1 vccd1 vccd1 _5091_/X sky130_fd_sc_hd__or4_1
XFILLER_37_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8850_ _8850_/A _4363_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[29] sky130_fd_sc_hd__ebufn_8
X_7801_ _7801_/A _7801_/B vssd1 vssd1 vccd1 vccd1 _7804_/A sky130_fd_sc_hd__xnor2_1
XFILLER_52_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5993_ _5993_/A _6259_/A vssd1 vssd1 vccd1 vccd1 _6000_/A sky130_fd_sc_hd__nor2_1
XFILLER_91_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7732_ _8205_/A _7886_/A vssd1 vssd1 vccd1 vccd1 _7760_/A sky130_fd_sc_hd__nand2_1
X_4944_ _5172_/C vssd1 vssd1 vccd1 vccd1 _5135_/C sky130_fd_sc_hd__clkbuf_2
X_7663_ _8057_/A _7671_/A _7666_/C vssd1 vssd1 vccd1 vccd1 _7665_/A sky130_fd_sc_hd__a21oi_1
X_4875_ _5104_/B _5006_/A vssd1 vssd1 vccd1 vccd1 _4959_/A sky130_fd_sc_hd__or2_1
X_6614_ _6656_/B vssd1 vssd1 vccd1 vccd1 _6614_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7594_ _7594_/A _7594_/B vssd1 vssd1 vccd1 vccd1 _7596_/A sky130_fd_sc_hd__nor2_1
X_6545_ _6545_/A _6545_/B vssd1 vssd1 vccd1 vccd1 _6545_/X sky130_fd_sc_hd__or2_1
X_8215_ _8132_/A _8212_/B _8131_/B _8214_/Y vssd1 vssd1 vccd1 vccd1 _8238_/A sky130_fd_sc_hd__o31ai_4
X_6476_ _8637_/Q _8636_/Q _8644_/Q vssd1 vssd1 vccd1 vccd1 _6477_/C sky130_fd_sc_hd__or3_1
X_5427_ _5421_/A _5419_/X _5426_/Y _5296_/X vssd1 vssd1 vccd1 vccd1 _8649_/D sky130_fd_sc_hd__o211a_1
X_8146_ _8363_/A _8146_/B vssd1 vssd1 vccd1 vccd1 _8151_/A sky130_fd_sc_hd__xor2_1
X_5358_ _8637_/Q _5360_/C _5357_/X vssd1 vssd1 vccd1 vccd1 _5359_/B sky130_fd_sc_hd__o21ai_1
XFILLER_101_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8077_ _8141_/A vssd1 vssd1 vccd1 vccd1 _8147_/A sky130_fd_sc_hd__clkbuf_2
XINSDIODE2_3 _5017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7028_ _7092_/A _7174_/B vssd1 vssd1 vccd1 vccd1 _7114_/B sky130_fd_sc_hd__nor2_2
X_5289_ _8717_/Q _5285_/X _5288_/X _5283_/X vssd1 vssd1 vccd1 vccd1 _8618_/D sky130_fd_sc_hd__o211a_1
XFILLER_28_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8814__92 vssd1 vssd1 vccd1 vccd1 _8814__92/HI _8923_/A sky130_fd_sc_hd__conb_1
XFILLER_74_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4660_ _4781_/A _4660_/B _4930_/A _4782_/A vssd1 vssd1 vccd1 vccd1 _4739_/A sky130_fd_sc_hd__or4b_2
X_4591_ _4598_/C _4646_/A _4591_/C vssd1 vssd1 vccd1 vccd1 _4592_/A sky130_fd_sc_hd__and3b_1
X_6330_ _6325_/X _6329_/X _4743_/X _8654_/Q vssd1 vssd1 vccd1 vccd1 _8654_/D sky130_fd_sc_hd__o2bb2a_1
XFILLER_6_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6261_ _6261_/A _6261_/B vssd1 vssd1 vccd1 vccd1 _6262_/B sky130_fd_sc_hd__xnor2_1
XFILLER_88_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8000_ _8074_/A _8000_/B vssd1 vssd1 vccd1 vccd1 _8001_/C sky130_fd_sc_hd__xor2_1
X_6192_ _6192_/A _6192_/B vssd1 vssd1 vccd1 vccd1 _6193_/B sky130_fd_sc_hd__xor2_1
X_5212_ _5129_/X _5210_/X _5212_/S vssd1 vssd1 vccd1 vccd1 _5213_/C sky130_fd_sc_hd__mux2_1
XFILLER_69_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5143_ _5143_/A _5143_/B vssd1 vssd1 vccd1 vccd1 _5144_/B sky130_fd_sc_hd__nor2_1
XFILLER_96_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5074_ _5214_/B _5074_/B _5149_/B _5193_/C vssd1 vssd1 vccd1 vccd1 _5074_/X sky130_fd_sc_hd__or4_1
X_8902_ _8902_/A _4420_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[11] sky130_fd_sc_hd__ebufn_8
XFILLER_37_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8833_ _8833_/A _4343_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[12] sky130_fd_sc_hd__ebufn_8
XFILLER_25_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5976_ _5976_/A _5976_/B vssd1 vssd1 vccd1 vccd1 _6025_/A sky130_fd_sc_hd__xor2_1
XFILLER_40_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7715_ _7745_/A _7745_/B vssd1 vssd1 vccd1 vccd1 _7884_/A sky130_fd_sc_hd__xnor2_2
X_8695_ input3/X _8695_/D vssd1 vssd1 vccd1 vccd1 _8695_/Q sky130_fd_sc_hd__dfxtp_1
X_4927_ _5115_/B _4939_/A vssd1 vssd1 vccd1 vccd1 _4928_/B sky130_fd_sc_hd__nor2_1
XFILLER_40_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7646_ _7664_/A _7682_/A vssd1 vssd1 vccd1 vccd1 _7816_/A sky130_fd_sc_hd__nor2_2
X_4858_ _5202_/A _5116_/B vssd1 vssd1 vccd1 vccd1 _5120_/A sky130_fd_sc_hd__or2_1
XFILLER_20_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7577_ _7658_/A _7552_/A _7576_/Y _7615_/B vssd1 vssd1 vccd1 vccd1 _7577_/X sky130_fd_sc_hd__a31o_1
X_4789_ _4789_/A _4822_/C vssd1 vssd1 vccd1 vccd1 _4848_/A sky130_fd_sc_hd__nor2_1
X_6528_ _6523_/A _6523_/B _6521_/B vssd1 vssd1 vccd1 vccd1 _6529_/B sky130_fd_sc_hd__a21oi_1
X_6459_ _8682_/Q _6459_/B _6459_/C vssd1 vssd1 vccd1 vccd1 _6463_/B sky130_fd_sc_hd__and3_1
X_8129_ _8225_/A _8130_/B vssd1 vssd1 vccd1 vccd1 _8212_/B sky130_fd_sc_hd__and2_2
XFILLER_102_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5830_ _5956_/A _5983_/A _6180_/B _5829_/Y vssd1 vssd1 vccd1 vccd1 _5831_/B sky130_fd_sc_hd__o31a_1
XFILLER_61_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5761_ _5954_/B _6284_/S _5777_/B vssd1 vssd1 vccd1 vccd1 _5764_/A sky130_fd_sc_hd__o21a_1
XFILLER_22_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8480_ _8480_/A _8480_/B vssd1 vssd1 vccd1 vccd1 _8481_/B sky130_fd_sc_hd__xnor2_1
X_7500_ _7505_/A _7505_/C vssd1 vssd1 vccd1 vccd1 _7501_/B sky130_fd_sc_hd__xnor2_1
X_4712_ _4716_/B _4712_/B _4712_/C vssd1 vssd1 vccd1 vccd1 _4713_/A sky130_fd_sc_hd__and3b_1
X_7431_ _7431_/A _7431_/B vssd1 vssd1 vccd1 vccd1 _7436_/A sky130_fd_sc_hd__xor2_1
X_5692_ _6107_/B _5692_/B vssd1 vssd1 vccd1 vccd1 _6046_/B sky130_fd_sc_hd__xnor2_2
X_4643_ _4645_/B _4643_/B vssd1 vssd1 vccd1 vccd1 _8589_/D sky130_fd_sc_hd__nor2_1
X_7362_ _7362_/A _7362_/B vssd1 vssd1 vccd1 vccd1 _7363_/B sky130_fd_sc_hd__xor2_1
X_4574_ _8572_/Q _8571_/Q vssd1 vssd1 vccd1 vccd1 _4587_/A sky130_fd_sc_hd__or2_1
X_7293_ _7293_/A _7293_/B vssd1 vssd1 vccd1 vccd1 _7294_/B sky130_fd_sc_hd__nand2_1
X_6313_ _6316_/A _6316_/B _6164_/X vssd1 vssd1 vccd1 vccd1 _6314_/B sky130_fd_sc_hd__a21o_1
X_6244_ _6244_/A _6244_/B vssd1 vssd1 vccd1 vccd1 _6244_/Y sky130_fd_sc_hd__nand2_1
XFILLER_97_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6175_ _6024_/A _6175_/B vssd1 vssd1 vccd1 vccd1 _6175_/X sky130_fd_sc_hd__and2b_1
XFILLER_97_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5126_ _5100_/X _5113_/Y _5125_/X _5060_/A vssd1 vssd1 vccd1 vccd1 _5126_/X sky130_fd_sc_hd__a31o_1
XFILLER_84_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5057_ _5057_/A _5229_/D _5057_/C _5057_/D vssd1 vssd1 vccd1 vccd1 _5058_/B sky130_fd_sc_hd__or4_1
XFILLER_72_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5959_ _5959_/A _6183_/A vssd1 vssd1 vccd1 vccd1 _5968_/B sky130_fd_sc_hd__xor2_1
XFILLER_21_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8678_ input3/X _8678_/D vssd1 vssd1 vccd1 vccd1 _8678_/Q sky130_fd_sc_hd__dfxtp_1
X_7629_ _8605_/Q _8708_/Q vssd1 vssd1 vccd1 vccd1 _7649_/A sky130_fd_sc_hd__nand2b_2
XFILLER_96_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7980_ _7980_/A _8021_/A _7980_/C vssd1 vssd1 vccd1 vccd1 _8021_/B sky130_fd_sc_hd__nand3_1
XFILLER_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6931_ _6931_/A _6931_/B vssd1 vssd1 vccd1 vccd1 _6932_/C sky130_fd_sc_hd__xor2_1
XFILLER_81_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6862_ _6862_/A vssd1 vssd1 vccd1 vccd1 _6880_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_34_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8601_ input3/X _8601_/D vssd1 vssd1 vccd1 vccd1 _8601_/Q sky130_fd_sc_hd__dfxtp_2
X_5813_ _5887_/B _5813_/B vssd1 vssd1 vccd1 vccd1 _5814_/B sky130_fd_sc_hd__or2_1
X_8532_ _8533_/A _8533_/B vssd1 vssd1 vccd1 vccd1 _8532_/Y sky130_fd_sc_hd__nor2_1
X_6793_ _7046_/A vssd1 vssd1 vccd1 vccd1 _7378_/B sky130_fd_sc_hd__clkbuf_2
X_5744_ _5744_/A _5744_/B vssd1 vssd1 vccd1 vccd1 _5786_/B sky130_fd_sc_hd__xor2_2
X_8463_ _8462_/B _8462_/C _8462_/Y vssd1 vssd1 vccd1 vccd1 _8464_/B sky130_fd_sc_hd__a21oi_1
X_5675_ _5675_/A _5675_/B vssd1 vssd1 vccd1 vccd1 _5746_/B sky130_fd_sc_hd__xor2_1
X_8394_ _8118_/A _7727_/X _8462_/A vssd1 vssd1 vccd1 vccd1 _8397_/A sky130_fd_sc_hd__a21oi_1
X_7414_ _7452_/A _7452_/B vssd1 vssd1 vccd1 vccd1 _7482_/A sky130_fd_sc_hd__xnor2_1
X_4626_ _8584_/Q _4628_/C _4646_/A vssd1 vssd1 vccd1 vccd1 _4626_/Y sky130_fd_sc_hd__o21ai_1
X_7345_ _7345_/A _7345_/B _7345_/C vssd1 vssd1 vccd1 vccd1 _7345_/X sky130_fd_sc_hd__or3_1
X_4557_ _8622_/Q _4563_/B vssd1 vssd1 vccd1 vccd1 _4558_/A sky130_fd_sc_hd__and2_1
XFILLER_1_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7276_ _7276_/A _7276_/B vssd1 vssd1 vccd1 vccd1 _7276_/Y sky130_fd_sc_hd__nor2_1
X_4488_ _8608_/Q vssd1 vssd1 vccd1 vccd1 _6617_/A sky130_fd_sc_hd__buf_2
XFILLER_103_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6227_ _5587_/Y _6226_/Y _6227_/S vssd1 vssd1 vccd1 vccd1 _6228_/B sky130_fd_sc_hd__mux2_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6158_ _6163_/A _6164_/D vssd1 vssd1 vccd1 vccd1 _6159_/B sky130_fd_sc_hd__xor2_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5109_ _5194_/A _5109_/B vssd1 vssd1 vccd1 vccd1 _5110_/D sky130_fd_sc_hd__or2_1
XFILLER_85_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6089_ _6134_/A _6134_/B vssd1 vssd1 vccd1 vccd1 _6135_/A sky130_fd_sc_hd__nor2_1
XFILLER_72_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8775__53 vssd1 vssd1 vccd1 vccd1 _8775__53/HI _8884_/A sky130_fd_sc_hd__conb_1
XFILLER_44_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5460_ _5460_/A _5460_/B vssd1 vssd1 vccd1 vccd1 _5486_/A sky130_fd_sc_hd__nor2_4
X_4411_ _4414_/A vssd1 vssd1 vccd1 vccd1 _4411_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5391_ _5391_/A vssd1 vssd1 vccd1 vccd1 _8645_/D sky130_fd_sc_hd__clkinv_2
X_7130_ _7042_/A _7042_/B _7129_/X vssd1 vssd1 vccd1 vccd1 _7131_/B sky130_fd_sc_hd__a21o_1
X_4342_ _4346_/A vssd1 vssd1 vccd1 vccd1 _4342_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7061_ _7060_/A _7060_/C _7060_/B vssd1 vssd1 vccd1 vccd1 _7063_/B sky130_fd_sc_hd__a21o_1
XFILLER_98_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6012_ _6011_/B _6012_/B vssd1 vssd1 vccd1 vccd1 _6013_/B sky130_fd_sc_hd__and2b_1
.ends

