* NGSPICE file created from wrapped_vgademo_on_fpga.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_8 abstract view
.subckt sky130_fd_sc_hd__ebufn_8 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_1 abstract view
.subckt sky130_fd_sc_hd__o311ai_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_4 abstract view
.subckt sky130_fd_sc_hd__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_4 abstract view
.subckt sky130_fd_sc_hd__nor2b_4 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_1 abstract view
.subckt sky130_fd_sc_hd__nor2b_1 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_2 abstract view
.subckt sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

.subckt wrapped_vgademo_on_fpga active io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21]
+ io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29]
+ io_in[2] io_in[30] io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37]
+ io_in[3] io_in[4] io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10]
+ io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18]
+ io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25]
+ io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32]
+ io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5]
+ io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12]
+ io_out[13] io_out[14] io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1]
+ io_out[20] io_out[21] io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27]
+ io_out[28] io_out[29] io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34]
+ io_out[35] io_out[36] io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ io_out[8] io_out[9] la1_data_in[0] la1_data_in[10] la1_data_in[11] la1_data_in[12]
+ la1_data_in[13] la1_data_in[14] la1_data_in[15] la1_data_in[16] la1_data_in[17]
+ la1_data_in[18] la1_data_in[19] la1_data_in[1] la1_data_in[20] la1_data_in[21] la1_data_in[22]
+ la1_data_in[23] la1_data_in[24] la1_data_in[25] la1_data_in[26] la1_data_in[27]
+ la1_data_in[28] la1_data_in[29] la1_data_in[2] la1_data_in[30] la1_data_in[31] la1_data_in[3]
+ la1_data_in[4] la1_data_in[5] la1_data_in[6] la1_data_in[7] la1_data_in[8] la1_data_in[9]
+ la1_data_out[0] la1_data_out[10] la1_data_out[11] la1_data_out[12] la1_data_out[13]
+ la1_data_out[14] la1_data_out[15] la1_data_out[16] la1_data_out[17] la1_data_out[18]
+ la1_data_out[19] la1_data_out[1] la1_data_out[20] la1_data_out[21] la1_data_out[22]
+ la1_data_out[23] la1_data_out[24] la1_data_out[25] la1_data_out[26] la1_data_out[27]
+ la1_data_out[28] la1_data_out[29] la1_data_out[2] la1_data_out[30] la1_data_out[31]
+ la1_data_out[3] la1_data_out[4] la1_data_out[5] la1_data_out[6] la1_data_out[7]
+ la1_data_out[8] la1_data_out[9] la1_oenb[0] la1_oenb[10] la1_oenb[11] la1_oenb[12]
+ la1_oenb[13] la1_oenb[14] la1_oenb[15] la1_oenb[16] la1_oenb[17] la1_oenb[18] la1_oenb[19]
+ la1_oenb[1] la1_oenb[20] la1_oenb[21] la1_oenb[22] la1_oenb[23] la1_oenb[24] la1_oenb[25]
+ la1_oenb[26] la1_oenb[27] la1_oenb[28] la1_oenb[29] la1_oenb[2] la1_oenb[30] la1_oenb[31]
+ la1_oenb[3] la1_oenb[4] la1_oenb[5] la1_oenb[6] la1_oenb[7] la1_oenb[8] la1_oenb[9]
+ vccd1 vssd1 wb_clk_i
XTAP_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7963_ _8064_/A _7963_/B vssd1 vssd1 vccd1 vccd1 _7964_/B sky130_fd_sc_hd__xor2_1
X_6914_ _6914_/A _6914_/B _6914_/C vssd1 vssd1 vccd1 vccd1 _6916_/B sky130_fd_sc_hd__and3_1
XFILLER_54_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7894_ _7942_/A _7942_/B vssd1 vssd1 vccd1 vccd1 _7903_/A sky130_fd_sc_hd__xnor2_4
XFILLER_23_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6845_ _6893_/A _6846_/B vssd1 vssd1 vccd1 vccd1 _6854_/A sky130_fd_sc_hd__nand2_1
X_6776_ _7079_/A vssd1 vssd1 vccd1 vccd1 _7310_/S sky130_fd_sc_hd__clkbuf_2
X_8515_ input3/X _8515_/D vssd1 vssd1 vccd1 vccd1 _8515_/Q sky130_fd_sc_hd__dfxtp_1
X_5727_ _5765_/A _5727_/B vssd1 vssd1 vccd1 vccd1 _5758_/B sky130_fd_sc_hd__xnor2_1
X_8446_ input3/X _8446_/D vssd1 vssd1 vccd1 vccd1 _8446_/Q sky130_fd_sc_hd__dfxtp_1
X_5658_ _5659_/A _5659_/B vssd1 vssd1 vccd1 vccd1 _6053_/B sky130_fd_sc_hd__nor2_1
X_4609_ _4609_/A vssd1 vssd1 vccd1 vccd1 _4619_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_8377_ _8381_/B _8377_/B vssd1 vssd1 vccd1 vccd1 _8378_/D sky130_fd_sc_hd__or2_1
X_5589_ _6082_/A _5590_/A vssd1 vssd1 vccd1 vccd1 _6249_/A sky130_fd_sc_hd__xor2_1
XFILLER_89_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7328_ _7328_/A _7328_/B vssd1 vssd1 vccd1 vccd1 _7329_/B sky130_fd_sc_hd__xor2_1
X_7259_ _7259_/A _7259_/B vssd1 vssd1 vccd1 vccd1 _7343_/A sky130_fd_sc_hd__nor2_1
XFILLER_77_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4960_ _4960_/A _4968_/A _5031_/C vssd1 vssd1 vccd1 vccd1 _5025_/A sky130_fd_sc_hd__or3_1
X_4891_ _5088_/A _5171_/B _4891_/C _5164_/B vssd1 vssd1 vccd1 vccd1 _4891_/X sky130_fd_sc_hd__or4_1
XFILLER_17_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6630_ _6627_/A _6627_/B _6627_/C _6606_/A _6539_/A vssd1 vssd1 vccd1 vccd1 _6736_/A
+ sky130_fd_sc_hd__a311o_1
X_6561_ _6999_/A _6999_/B _6479_/A vssd1 vssd1 vccd1 vccd1 _6652_/A sky130_fd_sc_hd__a21o_1
X_8300_ _8300_/A _8300_/B vssd1 vssd1 vccd1 vccd1 _8352_/A sky130_fd_sc_hd__xnor2_2
X_5512_ _6025_/A vssd1 vssd1 vccd1 vccd1 _5940_/A sky130_fd_sc_hd__buf_2
X_6492_ _7180_/A vssd1 vssd1 vccd1 vccd1 _7233_/A sky130_fd_sc_hd__buf_2
X_8231_ _8231_/A _8231_/B vssd1 vssd1 vccd1 vccd1 _8233_/C sky130_fd_sc_hd__xor2_1
X_5443_ _6281_/A _7575_/B _5459_/A _5459_/B _5437_/A vssd1 vssd1 vccd1 vccd1 _5444_/B
+ sky130_fd_sc_hd__a221o_1
X_8162_ _8282_/A _8282_/B vssd1 vssd1 vccd1 vccd1 _8163_/B sky130_fd_sc_hd__xnor2_1
X_5374_ _5374_/A _7494_/B vssd1 vssd1 vccd1 vccd1 _5417_/B sky130_fd_sc_hd__nand2_1
X_4325_ _4326_/A vssd1 vssd1 vccd1 vccd1 _4325_/Y sky130_fd_sc_hd__inv_2
X_7113_ _7156_/A _7156_/B _7112_/X vssd1 vssd1 vccd1 vccd1 _7134_/A sky130_fd_sc_hd__o21a_1
X_8093_ _8299_/A _8093_/B vssd1 vssd1 vccd1 vccd1 _8093_/Y sky130_fd_sc_hd__nor2_1
XFILLER_86_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7044_ _7044_/A _7044_/B vssd1 vssd1 vccd1 vccd1 _7045_/B sky130_fd_sc_hd__and2_1
XFILLER_47_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7946_ _7962_/A _7950_/A vssd1 vssd1 vccd1 vccd1 _8063_/B sky130_fd_sc_hd__or2_2
X_7877_ _7878_/B _7877_/B vssd1 vssd1 vccd1 vccd1 _7877_/X sky130_fd_sc_hd__and2b_1
X_6828_ _6828_/A _6828_/B vssd1 vssd1 vccd1 vccd1 _6873_/A sky130_fd_sc_hd__xnor2_2
XFILLER_23_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6759_ _6879_/B _6879_/C _6879_/A vssd1 vssd1 vccd1 vccd1 _6773_/A sky130_fd_sc_hd__a21bo_1
XFILLER_10_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8429_ _8424_/A _8428_/X _8429_/S vssd1 vssd1 vccd1 vccd1 _8430_/B sky130_fd_sc_hd__mux2_1
XFILLER_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5090_ _5090_/A _5090_/B _5117_/B vssd1 vssd1 vccd1 vccd1 _5118_/B sky130_fd_sc_hd__or3_1
XFILLER_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8780_ _8780_/A _4374_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[27] sky130_fd_sc_hd__ebufn_8
X_7800_ _8206_/B _7800_/B vssd1 vssd1 vccd1 vccd1 _8372_/B sky130_fd_sc_hd__xnor2_1
X_5992_ _5992_/A _5992_/B vssd1 vssd1 vccd1 vccd1 _5993_/B sky130_fd_sc_hd__xnor2_2
XFILLER_37_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4943_ _5088_/A _4943_/B vssd1 vssd1 vccd1 vccd1 _4947_/C sky130_fd_sc_hd__or2_1
XFILLER_52_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7731_ _7731_/A _7844_/A vssd1 vssd1 vccd1 vccd1 _7734_/A sky130_fd_sc_hd__nor2_1
X_7662_ _7769_/A _7712_/C vssd1 vssd1 vccd1 vccd1 _7664_/B sky130_fd_sc_hd__xnor2_1
X_4874_ _4839_/A _4869_/B _5112_/B _4868_/X _4873_/X vssd1 vssd1 vccd1 vccd1 _4874_/X
+ sky130_fd_sc_hd__o41a_1
X_6613_ _6640_/A _6622_/B _7032_/C _7039_/B vssd1 vssd1 vccd1 vccd1 _6616_/B sky130_fd_sc_hd__o31ai_2
X_7593_ _7899_/A _7952_/A _7954_/A vssd1 vssd1 vccd1 vccd1 _7717_/B sky130_fd_sc_hd__o21ai_1
X_6544_ _8553_/Q vssd1 vssd1 vccd1 vccd1 _6603_/A sky130_fd_sc_hd__inv_2
X_6475_ _8562_/Q _7559_/B vssd1 vssd1 vccd1 vccd1 _6475_/X sky130_fd_sc_hd__and2b_1
XFILLER_9_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8214_ _8356_/A _8213_/X _8356_/B vssd1 vssd1 vccd1 vccd1 _8214_/X sky130_fd_sc_hd__o21ba_1
X_5426_ _5426_/A _5426_/B vssd1 vssd1 vccd1 vccd1 _5427_/B sky130_fd_sc_hd__xnor2_1
XFILLER_59_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5357_ _5362_/A _5357_/B _5357_/C vssd1 vssd1 vccd1 vccd1 _5367_/S sky130_fd_sc_hd__nand3_2
X_8145_ _7756_/B _8273_/A _7899_/X vssd1 vssd1 vccd1 vccd1 _8258_/A sky130_fd_sc_hd__o21a_1
X_4308_ _4308_/A vssd1 vssd1 vccd1 vccd1 _4308_/Y sky130_fd_sc_hd__inv_2
X_5288_ _5290_/B _5288_/B vssd1 vssd1 vccd1 vccd1 _8503_/D sky130_fd_sc_hd__nor2_1
XINSDIODE2_4 _7239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8076_ _8076_/A _8134_/B vssd1 vssd1 vccd1 vccd1 _8116_/B sky130_fd_sc_hd__xnor2_1
XFILLER_87_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7027_ _6961_/B _7024_/X _7023_/Y _7021_/Y vssd1 vssd1 vccd1 vccd1 _7028_/C sky130_fd_sc_hd__a211o_1
X_8672__88 vssd1 vssd1 vccd1 vccd1 _8672__88/HI _8781_/A sky130_fd_sc_hd__conb_1
XFILLER_28_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7929_ _7930_/A _7930_/C _7930_/B vssd1 vssd1 vccd1 vccd1 _7993_/A sky130_fd_sc_hd__a21o_1
XFILLER_43_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4590_ _4735_/B _4882_/A _4675_/B vssd1 vssd1 vccd1 vccd1 _4747_/A sky130_fd_sc_hd__or3_2
XFILLER_9_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6260_ _6263_/S _6259_/Y _6264_/A _6264_/B _6264_/C vssd1 vssd1 vccd1 vccd1 _6260_/X
+ sky130_fd_sc_hd__a2111o_1
X_5211_ _8557_/Q _5202_/X _5210_/X _5200_/X vssd1 vssd1 vccd1 vccd1 _8482_/D sky130_fd_sc_hd__o211a_1
X_6191_ _5846_/A _5932_/B _6189_/Y _6190_/Y vssd1 vssd1 vccd1 vccd1 _6192_/B sky130_fd_sc_hd__o31a_1
XFILLER_96_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5142_ _5153_/A _5151_/B _5162_/B vssd1 vssd1 vccd1 vccd1 _5142_/X sky130_fd_sc_hd__or3_1
XFILLER_96_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5073_ _5073_/A vssd1 vssd1 vccd1 vccd1 _5073_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8763_ _8763_/A _4349_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[10] sky130_fd_sc_hd__ebufn_8
X_5975_ _5976_/A _6126_/B vssd1 vssd1 vccd1 vccd1 _5975_/X sky130_fd_sc_hd__and2_1
X_4926_ _5153_/A vssd1 vssd1 vccd1 vccd1 _5012_/A sky130_fd_sc_hd__clkbuf_2
X_8694_ _8694_/A _4273_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[11] sky130_fd_sc_hd__ebufn_8
X_7714_ _7715_/A _7715_/B vssd1 vssd1 vccd1 vccd1 _8207_/A sky130_fd_sc_hd__or2_1
X_4857_ _5132_/B _5132_/C _5148_/B _5149_/B vssd1 vssd1 vccd1 vccd1 _5135_/C sky130_fd_sc_hd__or4_1
XFILLER_20_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7645_ _7822_/A _7645_/B vssd1 vssd1 vccd1 vccd1 _7647_/A sky130_fd_sc_hd__nand2_2
XFILLER_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7576_ _7576_/A _7576_/B vssd1 vssd1 vccd1 vccd1 _7606_/A sky130_fd_sc_hd__nand2_1
X_4788_ _5010_/A _5138_/A vssd1 vssd1 vccd1 vccd1 _4968_/A sky130_fd_sc_hd__or2_1
X_6527_ _6513_/X _6570_/B _6570_/C _6512_/A _6506_/A vssd1 vssd1 vccd1 vccd1 _6557_/A
+ sky130_fd_sc_hd__a311o_1
XFILLER_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6458_ _6541_/A _8549_/Q vssd1 vssd1 vccd1 vccd1 _6459_/D sky130_fd_sc_hd__or2_1
XFILLER_79_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6389_ _6387_/Y _6389_/B vssd1 vssd1 vccd1 vccd1 _6390_/A sky130_fd_sc_hd__and2b_1
X_5409_ _5538_/A _5537_/B vssd1 vssd1 vccd1 vccd1 _5565_/A sky130_fd_sc_hd__or2_1
XFILLER_87_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8128_ _8257_/A _8128_/B vssd1 vssd1 vccd1 vccd1 _8129_/B sky130_fd_sc_hd__or2_1
XFILLER_85_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8059_ _7958_/X _7967_/B _7959_/A vssd1 vssd1 vccd1 vccd1 _8075_/A sky130_fd_sc_hd__a21oi_1
XFILLER_18_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5760_ _5824_/A vssd1 vssd1 vccd1 vccd1 _6021_/A sky130_fd_sc_hd__buf_2
X_4711_ _4711_/A _4711_/B vssd1 vssd1 vccd1 vccd1 _5131_/B sky130_fd_sc_hd__or2_1
XFILLER_61_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5691_ _6053_/A _5691_/B _5711_/B vssd1 vssd1 vccd1 vccd1 _5692_/B sky130_fd_sc_hd__or3_1
X_4642_ _4642_/A _4862_/B vssd1 vssd1 vccd1 vccd1 _4711_/B sky130_fd_sc_hd__nand2_1
X_7430_ _8423_/A _8428_/A _7428_/X _7429_/X _4510_/A vssd1 vssd1 vccd1 vccd1 _8568_/D
+ sky130_fd_sc_hd__o311ai_1
X_7361_ _7352_/X _7360_/Y _7354_/Y _7350_/Y vssd1 vssd1 vccd1 vccd1 _7361_/X sky130_fd_sc_hd__o211a_1
X_4573_ _8452_/Q _4574_/B vssd1 vssd1 vccd1 vccd1 _4575_/B sky130_fd_sc_hd__or2_1
X_6312_ _8539_/Q _6310_/X _6371_/B vssd1 vssd1 vccd1 vccd1 _6312_/X sky130_fd_sc_hd__a21o_1
X_7292_ _6622_/B _6980_/A _7292_/S vssd1 vssd1 vccd1 vccd1 _7293_/B sky130_fd_sc_hd__mux2_1
X_6243_ _6243_/A _6243_/B vssd1 vssd1 vccd1 vccd1 _6243_/Y sky130_fd_sc_hd__nand2_1
XFILLER_69_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6174_ _6174_/A _6174_/B vssd1 vssd1 vccd1 vccd1 _6174_/Y sky130_fd_sc_hd__nor2_1
X_5125_ _5125_/A _5135_/B _5125_/C vssd1 vssd1 vccd1 vccd1 _5125_/X sky130_fd_sc_hd__or3_1
XFILLER_57_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5056_ _5064_/B _5149_/B _5056_/C vssd1 vssd1 vccd1 vccd1 _5057_/B sky130_fd_sc_hd__or3_1
XFILLER_57_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8642__58 vssd1 vssd1 vccd1 vccd1 _8642__58/HI _8751_/A sky130_fd_sc_hd__conb_1
XFILLER_84_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8746_ _8746_/A _4336_/Y vssd1 vssd1 vccd1 vccd1 io_out[31] sky130_fd_sc_hd__ebufn_8
X_5958_ _5967_/A _5967_/B vssd1 vssd1 vccd1 vccd1 _5959_/B sky130_fd_sc_hd__xor2_1
XFILLER_25_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4909_ _4909_/A _4909_/B _4771_/X vssd1 vssd1 vccd1 vccd1 _4975_/C sky130_fd_sc_hd__or3b_2
XFILLER_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5889_ _5889_/A _5889_/B vssd1 vssd1 vccd1 vccd1 _5890_/B sky130_fd_sc_hd__xor2_1
X_7628_ _8147_/A _8146_/A _8146_/B vssd1 vssd1 vccd1 vccd1 _8070_/A sky130_fd_sc_hd__or3_2
XFILLER_4_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7559_ _8582_/Q _7559_/B vssd1 vssd1 vccd1 vccd1 _7559_/X sky130_fd_sc_hd__and2b_1
XFILLER_20_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6930_ _6930_/A _6930_/B vssd1 vssd1 vccd1 vccd1 _6949_/B sky130_fd_sc_hd__and2_1
XFILLER_66_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6861_ _7282_/A _7282_/B vssd1 vssd1 vccd1 vccd1 _6862_/B sky130_fd_sc_hd__xor2_2
XFILLER_19_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6792_ _7310_/S _6792_/B _6792_/C vssd1 vssd1 vccd1 vccd1 _6794_/A sky130_fd_sc_hd__and3_1
XFILLER_62_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5812_ _5812_/A _5812_/B vssd1 vssd1 vccd1 vccd1 _5813_/B sky130_fd_sc_hd__nand2_1
XFILLER_62_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8531_ input3/X _8531_/D vssd1 vssd1 vccd1 vccd1 _8531_/Q sky130_fd_sc_hd__dfxtp_1
X_5743_ _5743_/A _5743_/B vssd1 vssd1 vccd1 vccd1 _5751_/B sky130_fd_sc_hd__xnor2_1
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8462_ input3/X _8462_/D vssd1 vssd1 vccd1 vccd1 _8462_/Q sky130_fd_sc_hd__dfxtp_4
X_5674_ _5673_/B _5673_/C _5673_/A vssd1 vssd1 vccd1 vccd1 _5676_/B sky130_fd_sc_hd__o21ai_1
XFILLER_30_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4625_ _6482_/B vssd1 vssd1 vccd1 vccd1 _4626_/A sky130_fd_sc_hd__inv_2
X_7413_ _7413_/A vssd1 vssd1 vccd1 vccd1 _8567_/D sky130_fd_sc_hd__clkbuf_1
X_8393_ _8581_/Q _8393_/B vssd1 vssd1 vccd1 vccd1 _8393_/Y sky130_fd_sc_hd__xnor2_1
X_7344_ _7344_/A _7344_/B vssd1 vssd1 vccd1 vccd1 _7344_/X sky130_fd_sc_hd__xor2_1
X_4556_ _8446_/Q _4557_/C _4555_/Y vssd1 vssd1 vccd1 vccd1 _8446_/D sky130_fd_sc_hd__a21oi_1
X_4487_ _8485_/Q _4491_/B vssd1 vssd1 vccd1 vccd1 _4488_/A sky130_fd_sc_hd__and2_1
XFILLER_89_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7275_ _6962_/A _6962_/B _6963_/B _7093_/A vssd1 vssd1 vccd1 vccd1 _7336_/A sky130_fd_sc_hd__o22a_1
XFILLER_89_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6226_ _6226_/A _6226_/B vssd1 vssd1 vccd1 vccd1 _6227_/B sky130_fd_sc_hd__xnor2_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6157_ _6195_/A _6195_/B vssd1 vssd1 vccd1 vccd1 _6158_/B sky130_fd_sc_hd__xnor2_1
X_5108_ _5179_/A _5030_/B _5103_/X _5107_/X vssd1 vssd1 vccd1 vccd1 _5109_/D sky130_fd_sc_hd__o31a_1
XFILLER_85_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6088_ _6088_/A _6088_/B vssd1 vssd1 vccd1 vccd1 _6233_/B sky130_fd_sc_hd__xor2_1
XFILLER_17_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5039_ _5138_/A _5039_/B vssd1 vssd1 vccd1 vccd1 _5117_/C sky130_fd_sc_hd__or2_1
XFILLER_72_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8729_ _8729_/A _4314_/Y vssd1 vssd1 vccd1 vccd1 io_out[14] sky130_fd_sc_hd__ebufn_8
XFILLER_9_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4410_ _4718_/A vssd1 vssd1 vccd1 vccd1 _4735_/A sky130_fd_sc_hd__clkbuf_1
X_5390_ _5686_/A _5800_/A vssd1 vssd1 vccd1 vccd1 _5426_/A sky130_fd_sc_hd__nand2_2
X_4341_ _4345_/A vssd1 vssd1 vccd1 vccd1 _4341_/Y sky130_fd_sc_hd__inv_2
X_7060_ _7060_/A _7060_/B vssd1 vssd1 vccd1 vccd1 _7114_/B sky130_fd_sc_hd__xor2_1
X_4272_ _4296_/A vssd1 vssd1 vccd1 vccd1 _4277_/A sky130_fd_sc_hd__clkbuf_2
X_6011_ _6011_/A _6011_/B vssd1 vssd1 vccd1 vccd1 _6044_/A sky130_fd_sc_hd__nand2_1
X_8612__28 vssd1 vssd1 vccd1 vccd1 _8612__28/HI _8707_/A sky130_fd_sc_hd__conb_1
XFILLER_27_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7962_ _7962_/A _8146_/A _8146_/B vssd1 vssd1 vccd1 vccd1 _7963_/B sky130_fd_sc_hd__or3_1
X_6913_ _6913_/A _6913_/B vssd1 vssd1 vccd1 vccd1 _6983_/A sky130_fd_sc_hd__xnor2_1
XFILLER_54_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7893_ _8142_/A _7893_/B vssd1 vssd1 vccd1 vccd1 _7942_/B sky130_fd_sc_hd__xnor2_2
XFILLER_23_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6844_ _6804_/A _7175_/B _6844_/S vssd1 vssd1 vccd1 vccd1 _6846_/B sky130_fd_sc_hd__mux2_1
XFILLER_52_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6775_ _6886_/A _6886_/B _6774_/X vssd1 vssd1 vccd1 vccd1 _6795_/A sky130_fd_sc_hd__o21a_1
XFILLER_22_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5726_ _5619_/A _5724_/Y _5725_/X vssd1 vssd1 vccd1 vccd1 _5727_/B sky130_fd_sc_hd__a21o_1
X_8514_ input3/X _8514_/D vssd1 vssd1 vccd1 vccd1 _8514_/Q sky130_fd_sc_hd__dfxtp_1
X_8445_ input3/X _8445_/D vssd1 vssd1 vccd1 vccd1 _8445_/Q sky130_fd_sc_hd__dfxtp_1
X_5657_ _5543_/A _5543_/B _5426_/A _5406_/B vssd1 vssd1 vccd1 vccd1 _5659_/B sky130_fd_sc_hd__o2bb2a_1
X_4608_ _5151_/A vssd1 vssd1 vccd1 vccd1 _4609_/A sky130_fd_sc_hd__clkbuf_2
X_8376_ _8375_/B _8376_/B vssd1 vssd1 vccd1 vccd1 _8377_/B sky130_fd_sc_hd__and2b_1
X_5588_ _6248_/A _5591_/B vssd1 vssd1 vccd1 vccd1 _5590_/A sky130_fd_sc_hd__nand2_1
X_7327_ _6647_/A _6647_/B _6560_/B _6714_/A vssd1 vssd1 vccd1 vccd1 _7328_/B sky130_fd_sc_hd__a22o_1
X_4539_ _8440_/Q _8441_/Q _4539_/C vssd1 vssd1 vccd1 vccd1 _4543_/B sky130_fd_sc_hd__and3_1
X_7258_ _7200_/B _7200_/C _7200_/A vssd1 vssd1 vccd1 vccd1 _7258_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_77_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6209_ _6209_/A _6209_/B vssd1 vssd1 vccd1 vccd1 _6210_/B sky130_fd_sc_hd__xnor2_1
X_7189_ _7191_/B _7191_/A vssd1 vssd1 vccd1 vccd1 _7196_/A sky130_fd_sc_hd__and2b_1
XFILLER_85_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8678__94 vssd1 vssd1 vccd1 vccd1 _8678__94/HI _8787_/A sky130_fd_sc_hd__conb_1
XFILLER_5_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4890_ _4890_/A vssd1 vssd1 vccd1 vccd1 _5164_/B sky130_fd_sc_hd__inv_2
X_6560_ _6647_/B _6560_/B vssd1 vssd1 vccd1 vccd1 _6702_/A sky130_fd_sc_hd__or2_1
X_5511_ _5609_/C vssd1 vssd1 vccd1 vccd1 _6025_/A sky130_fd_sc_hd__clkbuf_2
X_6491_ _7043_/A vssd1 vssd1 vccd1 vccd1 _7180_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_8_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8230_ _8306_/A _8305_/S vssd1 vssd1 vccd1 vccd1 _8233_/A sky130_fd_sc_hd__nor2_1
X_5442_ _5455_/A _5455_/B _5441_/X vssd1 vssd1 vccd1 vccd1 _5459_/B sky130_fd_sc_hd__a21o_2
X_8161_ _8074_/A _8074_/B _8160_/X vssd1 vssd1 vccd1 vccd1 _8282_/B sky130_fd_sc_hd__a21oi_1
X_5373_ _5373_/A vssd1 vssd1 vccd1 vccd1 _5417_/A sky130_fd_sc_hd__clkbuf_4
X_7112_ _7155_/A _7107_/B vssd1 vssd1 vccd1 vccd1 _7112_/X sky130_fd_sc_hd__or2b_1
X_4324_ _4326_/A vssd1 vssd1 vccd1 vccd1 _4324_/Y sky130_fd_sc_hd__inv_2
X_8092_ _8092_/A _8031_/B vssd1 vssd1 vccd1 vccd1 _8111_/B sky130_fd_sc_hd__or2b_1
XFILLER_86_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7043_ _7043_/A _7043_/B vssd1 vssd1 vccd1 vccd1 _7105_/A sky130_fd_sc_hd__nor2_2
XFILLER_86_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7945_ _7945_/A _7945_/B _7945_/C vssd1 vssd1 vccd1 vccd1 _7945_/X sky130_fd_sc_hd__or3_1
X_7876_ _7869_/A _7869_/B _7875_/X vssd1 vssd1 vccd1 vccd1 _7939_/A sky130_fd_sc_hd__a21o_1
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6827_ _6825_/Y _6827_/B vssd1 vssd1 vccd1 vccd1 _6828_/B sky130_fd_sc_hd__and2b_1
XFILLER_50_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6758_ _6758_/A _6816_/B _6758_/C vssd1 vssd1 vccd1 vccd1 _6879_/A sky130_fd_sc_hd__nand3_1
XFILLER_7_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6689_ _6690_/A _6690_/C _7294_/B vssd1 vssd1 vccd1 vccd1 _6791_/A sky130_fd_sc_hd__o21a_1
X_5709_ _5855_/A vssd1 vssd1 vccd1 vccd1 _5861_/A sky130_fd_sc_hd__clkinv_2
X_8428_ _8428_/A _8428_/B vssd1 vssd1 vccd1 vccd1 _8428_/X sky130_fd_sc_hd__or2_1
XFILLER_88_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8359_ _8359_/A _8359_/B _8359_/C vssd1 vssd1 vccd1 vccd1 _8362_/A sky130_fd_sc_hd__nand3_1
XFILLER_88_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5991_ _5989_/Y _5991_/B vssd1 vssd1 vccd1 vccd1 _5992_/B sky130_fd_sc_hd__and2b_1
XFILLER_24_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4942_ _4921_/X _4937_/X _4939_/X _4941_/X vssd1 vssd1 vccd1 vccd1 _4942_/X sky130_fd_sc_hd__o31a_1
X_7730_ _7742_/A _8147_/A vssd1 vssd1 vccd1 vccd1 _7860_/A sky130_fd_sc_hd__nor2_1
XFILLER_32_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7661_ _7783_/A _7661_/B vssd1 vssd1 vccd1 vccd1 _7712_/C sky130_fd_sc_hd__xnor2_1
X_4873_ _4873_/A _4969_/A _4955_/B _5136_/C vssd1 vssd1 vccd1 vccd1 _4873_/X sky130_fd_sc_hd__or4_1
XFILLER_60_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6612_ _6964_/C vssd1 vssd1 vccd1 vccd1 _7032_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_20_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7592_ _8317_/B _8054_/A vssd1 vssd1 vccd1 vccd1 _7954_/A sky130_fd_sc_hd__or2_1
XFILLER_20_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6543_ _8471_/Q _8554_/Q vssd1 vssd1 vccd1 vccd1 _6543_/X sky130_fd_sc_hd__or2b_1
X_6474_ _8562_/Q _7559_/B vssd1 vssd1 vccd1 vccd1 _6486_/B sky130_fd_sc_hd__xnor2_1
X_8213_ _8210_/A _8213_/B _8213_/C _8213_/D vssd1 vssd1 vccd1 vccd1 _8213_/X sky130_fd_sc_hd__and4b_1
X_5425_ _5648_/A _5855_/A vssd1 vssd1 vccd1 vccd1 _5426_/B sky130_fd_sc_hd__nor2_1
X_5356_ _5362_/A _5357_/B _5357_/C vssd1 vssd1 vccd1 vccd1 _5356_/X sky130_fd_sc_hd__a21o_1
X_8144_ _8248_/A _8248_/B vssd1 vssd1 vccd1 vccd1 _8163_/A sky130_fd_sc_hd__xnor2_1
X_4307_ _4308_/A vssd1 vssd1 vccd1 vccd1 _4307_/Y sky130_fd_sc_hd__inv_2
XINSDIODE2_5 _7244_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5287_ _8503_/Q _5286_/B _5230_/B vssd1 vssd1 vccd1 vccd1 _5288_/B sky130_fd_sc_hd__o21ai_1
X_8075_ _8075_/A _8133_/B vssd1 vssd1 vccd1 vccd1 _8134_/B sky130_fd_sc_hd__xnor2_1
X_7026_ _7026_/A vssd1 vssd1 vccd1 vccd1 _7146_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_74_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7928_ _8003_/A _7927_/X vssd1 vssd1 vccd1 vccd1 _7930_/B sky130_fd_sc_hd__or2b_1
XFILLER_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7859_ _7899_/A _8064_/A vssd1 vssd1 vccd1 vccd1 _7864_/A sky130_fd_sc_hd__nor2_1
XFILLER_23_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8648__64 vssd1 vssd1 vccd1 vccd1 _8648__64/HI _8757_/A sky130_fd_sc_hd__conb_1
XFILLER_93_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5210_ _8482_/Q _5217_/B vssd1 vssd1 vccd1 vccd1 _5210_/X sky130_fd_sc_hd__or2_1
X_6190_ _5930_/B _6189_/Y _5846_/Y vssd1 vssd1 vccd1 vccd1 _6190_/Y sky130_fd_sc_hd__o21bai_1
X_5141_ _4623_/X _4830_/Y _5121_/X _5140_/X _5175_/S vssd1 vssd1 vccd1 vccd1 _5141_/X
+ sky130_fd_sc_hd__o32a_1
X_5072_ _5072_/A _5109_/C _5093_/D vssd1 vssd1 vccd1 vccd1 _5073_/A sky130_fd_sc_hd__or3_1
XFILLER_96_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8762_ _8762_/A _4347_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[9] sky130_fd_sc_hd__ebufn_8
XFILLER_25_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5974_ _5581_/A _6243_/A _5984_/B vssd1 vssd1 vccd1 vccd1 _5983_/A sky130_fd_sc_hd__a21o_1
XFILLER_40_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7713_ _7710_/Y _7661_/B _7712_/X vssd1 vssd1 vccd1 vccd1 _7715_/B sky130_fd_sc_hd__a21oi_1
X_4925_ _5136_/A vssd1 vssd1 vccd1 vccd1 _5171_/A sky130_fd_sc_hd__clkbuf_2
X_8693_ _8693_/A _4270_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[10] sky130_fd_sc_hd__ebufn_8
X_4856_ _5030_/C vssd1 vssd1 vccd1 vccd1 _5149_/B sky130_fd_sc_hd__clkbuf_2
X_7644_ _7766_/A _7644_/B vssd1 vssd1 vccd1 vccd1 _7645_/B sky130_fd_sc_hd__nand2_1
X_7575_ _8405_/A _7575_/B vssd1 vssd1 vccd1 vccd1 _7576_/B sky130_fd_sc_hd__nand2_1
X_4787_ _5162_/B _4956_/C vssd1 vssd1 vccd1 vccd1 _5010_/A sky130_fd_sc_hd__or2_1
X_6526_ _6558_/A vssd1 vssd1 vccd1 vccd1 _7054_/A sky130_fd_sc_hd__buf_2
XFILLER_20_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6457_ _6541_/A _8549_/Q vssd1 vssd1 vccd1 vccd1 _6466_/B sky130_fd_sc_hd__nand2_1
X_6388_ _8546_/Q _6386_/A _6387_/Y _4668_/X vssd1 vssd1 vccd1 vccd1 _8546_/D sky130_fd_sc_hd__o211a_1
X_5408_ _5694_/A _5408_/B _5408_/C vssd1 vssd1 vccd1 vccd1 _5537_/B sky130_fd_sc_hd__and3_1
X_5339_ _8508_/Q _5339_/B vssd1 vssd1 vccd1 vccd1 _5341_/A sky130_fd_sc_hd__and2b_1
X_8127_ _8127_/A _8127_/B vssd1 vssd1 vccd1 vccd1 _8128_/B sky130_fd_sc_hd__and2_1
XFILLER_87_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8058_ _8129_/A _8058_/B vssd1 vssd1 vccd1 vccd1 _8076_/A sky130_fd_sc_hd__nand2_1
X_7009_ _7009_/A _7009_/B vssd1 vssd1 vccd1 vccd1 _7011_/B sky130_fd_sc_hd__xnor2_1
XFILLER_18_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4710_ _4711_/A _4711_/B vssd1 vssd1 vccd1 vccd1 _5131_/A sky130_fd_sc_hd__nand2_1
X_5690_ _6053_/A _5691_/B _5711_/B vssd1 vssd1 vccd1 vccd1 _5809_/A sky130_fd_sc_hd__o21ai_1
XFILLER_42_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4641_ _4638_/A _4640_/A _4640_/Y _4602_/X vssd1 vssd1 vccd1 vccd1 _8459_/D sky130_fd_sc_hd__o211a_1
XFILLER_30_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7360_ _7365_/B vssd1 vssd1 vccd1 vccd1 _7360_/Y sky130_fd_sc_hd__inv_2
X_4572_ _4574_/B _4572_/B vssd1 vssd1 vccd1 vccd1 _8451_/D sky130_fd_sc_hd__nor2_1
X_6311_ _8540_/Q vssd1 vssd1 vccd1 vccd1 _6371_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_7291_ _7291_/A _7291_/B vssd1 vssd1 vccd1 vccd1 _7292_/S sky130_fd_sc_hd__nor2_1
X_6242_ _6069_/X _6231_/Y _6240_/Y _6241_/X vssd1 vssd1 vccd1 vccd1 _6264_/C sky130_fd_sc_hd__a211o_2
X_6173_ _6167_/A _6173_/B vssd1 vssd1 vccd1 vccd1 _6173_/X sky130_fd_sc_hd__and2b_1
X_5124_ _5057_/B _5121_/X _5123_/X _4626_/A vssd1 vssd1 vccd1 vccd1 _5125_/C sky130_fd_sc_hd__o22a_1
XFILLER_69_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5055_ _5055_/A _5055_/B _5116_/B vssd1 vssd1 vccd1 vccd1 _5056_/C sky130_fd_sc_hd__or3_1
XFILLER_84_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8745_ _8745_/A _4335_/Y vssd1 vssd1 vccd1 vccd1 io_out[30] sky130_fd_sc_hd__ebufn_8
X_5957_ _5957_/A _5957_/B vssd1 vssd1 vccd1 vccd1 _5967_/B sky130_fd_sc_hd__xnor2_2
X_4908_ _4908_/A _4908_/B vssd1 vssd1 vccd1 vccd1 _4909_/A sky130_fd_sc_hd__and2_1
XFILLER_40_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5888_ _5888_/A _5888_/B vssd1 vssd1 vccd1 vccd1 _5889_/B sky130_fd_sc_hd__nand2_1
X_7627_ _7741_/A vssd1 vssd1 vccd1 vccd1 _8146_/B sky130_fd_sc_hd__clkbuf_2
X_4839_ _4839_/A _5089_/A vssd1 vssd1 vccd1 vccd1 _4839_/X sky130_fd_sc_hd__or2_1
X_7558_ _8582_/Q _7559_/B vssd1 vssd1 vccd1 vccd1 _7569_/B sky130_fd_sc_hd__xnor2_4
X_6509_ _6509_/A _6509_/B vssd1 vssd1 vccd1 vccd1 _7365_/A sky130_fd_sc_hd__xor2_2
X_7489_ _8426_/A _7489_/B vssd1 vssd1 vccd1 vccd1 _7489_/Y sky130_fd_sc_hd__nor2_1
XFILLER_96_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8618__34 vssd1 vssd1 vccd1 vccd1 _8618__34/HI _8713_/A sky130_fd_sc_hd__conb_1
XFILLER_88_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6860_ _6860_/A _7289_/B vssd1 vssd1 vccd1 vccd1 _7282_/B sky130_fd_sc_hd__xor2_2
X_6791_ _6791_/A _6791_/B _6789_/Y vssd1 vssd1 vccd1 vccd1 _6792_/C sky130_fd_sc_hd__or3b_1
XFILLER_62_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5811_ _5811_/A _5811_/B vssd1 vssd1 vccd1 vccd1 _5812_/A sky130_fd_sc_hd__nand2_1
XFILLER_22_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8530_ input3/X _8530_/D vssd1 vssd1 vccd1 vccd1 _8530_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5742_ _5754_/A _5754_/B vssd1 vssd1 vccd1 vccd1 _5743_/B sky130_fd_sc_hd__xnor2_1
X_8461_ input3/X _8461_/D vssd1 vssd1 vccd1 vccd1 _8461_/Q sky130_fd_sc_hd__dfxtp_2
X_5673_ _5673_/A _5673_/B _5673_/C vssd1 vssd1 vccd1 vccd1 _6070_/B sky130_fd_sc_hd__or3_1
X_4624_ _4624_/A _5016_/A vssd1 vssd1 vccd1 vccd1 _4862_/A sky130_fd_sc_hd__nor2_1
X_7412_ _7412_/A _7412_/B _7412_/C vssd1 vssd1 vccd1 vccd1 _7413_/A sky130_fd_sc_hd__and3_1
X_8392_ _8392_/A _8392_/B vssd1 vssd1 vccd1 vccd1 _8393_/B sky130_fd_sc_hd__nand2_1
X_7343_ _7343_/A _7217_/Y vssd1 vssd1 vccd1 vccd1 _7344_/A sky130_fd_sc_hd__or2b_1
X_4555_ _8446_/Q _4557_/C _4575_/A vssd1 vssd1 vccd1 vccd1 _4555_/Y sky130_fd_sc_hd__o21ai_1
X_4486_ _4486_/A vssd1 vssd1 vccd1 vccd1 _8738_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7274_ _7268_/A _7268_/B _7268_/C _7273_/Y vssd1 vssd1 vccd1 vccd1 _7337_/A sky130_fd_sc_hd__a31o_1
X_6225_ _6225_/A _6225_/B vssd1 vssd1 vccd1 vccd1 _6226_/B sky130_fd_sc_hd__nand2_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6156_ _6156_/A _6156_/B vssd1 vssd1 vccd1 vccd1 _6195_/B sky130_fd_sc_hd__xnor2_1
X_5107_ _5121_/A _5136_/B _5107_/C _5107_/D vssd1 vssd1 vccd1 vccd1 _5107_/X sky130_fd_sc_hd__or4_1
XFILLER_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6087_ _6087_/A _6090_/C vssd1 vssd1 vccd1 vccd1 _6233_/A sky130_fd_sc_hd__and2_1
X_5038_ _5012_/A _5091_/A _5037_/X _5028_/X vssd1 vssd1 vccd1 vccd1 _5038_/X sky130_fd_sc_hd__a211o_1
XFILLER_72_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8728_ _8728_/A _4313_/Y vssd1 vssd1 vccd1 vccd1 io_out[13] sky130_fd_sc_hd__ebufn_8
XFILLER_80_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6989_ _6989_/A _6989_/B vssd1 vssd1 vccd1 vccd1 _6992_/A sky130_fd_sc_hd__nor2_1
XFILLER_25_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4340_ _4358_/A vssd1 vssd1 vccd1 vccd1 _4345_/A sky130_fd_sc_hd__clkbuf_2
X_4271_ input1/X vssd1 vssd1 vccd1 vccd1 _4296_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_4_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6010_ _6010_/A _6010_/B vssd1 vssd1 vccd1 vccd1 _6011_/B sky130_fd_sc_hd__or2_1
XFILLER_79_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7961_ _7961_/A _8326_/B vssd1 vssd1 vccd1 vccd1 _7964_/A sky130_fd_sc_hd__nor2_1
XFILLER_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6912_ _6912_/A _6912_/B vssd1 vssd1 vccd1 vccd1 _6962_/A sky130_fd_sc_hd__xnor2_1
X_7892_ _7945_/B _7945_/C vssd1 vssd1 vccd1 vccd1 _7893_/B sky130_fd_sc_hd__nor2_1
X_6843_ _6971_/A vssd1 vssd1 vccd1 vccd1 _6893_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_62_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6774_ _6774_/A _6773_/A vssd1 vssd1 vccd1 vccd1 _6774_/X sky130_fd_sc_hd__or2b_1
X_8513_ input3/X _8513_/D vssd1 vssd1 vccd1 vccd1 _8513_/Q sky130_fd_sc_hd__dfxtp_1
X_5725_ _5764_/A _5825_/B _5825_/C _5724_/A _6025_/A vssd1 vssd1 vccd1 vccd1 _5725_/X
+ sky130_fd_sc_hd__o32a_1
X_5656_ _5699_/A _5699_/B vssd1 vssd1 vccd1 vccd1 _5662_/A sky130_fd_sc_hd__xnor2_1
X_8444_ input3/X _8444_/D vssd1 vssd1 vccd1 vccd1 _8444_/Q sky130_fd_sc_hd__dfxtp_1
X_4607_ _5102_/A vssd1 vssd1 vccd1 vccd1 _5151_/A sky130_fd_sc_hd__clkbuf_2
X_8375_ _8376_/B _8375_/B vssd1 vssd1 vccd1 vccd1 _8381_/B sky130_fd_sc_hd__and2b_1
X_5587_ _6247_/A _6247_/B vssd1 vssd1 vccd1 vccd1 _5591_/B sky130_fd_sc_hd__and2b_1
X_7326_ _6838_/A _6838_/B _7325_/X vssd1 vssd1 vccd1 vccd1 _7329_/A sky130_fd_sc_hd__a21oi_1
X_4538_ _8440_/Q _4539_/C _4537_/Y vssd1 vssd1 vccd1 vccd1 _8440_/D sky130_fd_sc_hd__a21oi_1
X_7257_ _7354_/A _7354_/B _7256_/Y vssd1 vssd1 vccd1 vccd1 _7344_/B sky130_fd_sc_hd__a21o_1
X_4469_ _4469_/A _4469_/B _4659_/A vssd1 vssd1 vccd1 vccd1 _4470_/D sky130_fd_sc_hd__and3_1
XFILLER_58_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6208_ _6208_/A _6208_/B vssd1 vssd1 vccd1 vccd1 _6209_/B sky130_fd_sc_hd__xnor2_1
X_7188_ _7177_/A _7177_/B _7177_/C _7211_/A vssd1 vssd1 vccd1 vccd1 _7191_/A sky130_fd_sc_hd__a31o_1
XFILLER_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6139_ _5518_/C _5829_/C _5930_/B vssd1 vssd1 vccd1 vccd1 _6198_/B sky130_fd_sc_hd__a21oi_1
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5510_ _5949_/A vssd1 vssd1 vccd1 vccd1 _5637_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6490_ _6584_/A vssd1 vssd1 vccd1 vccd1 _7043_/A sky130_fd_sc_hd__clkbuf_2
X_5441_ _8521_/Q _5441_/B vssd1 vssd1 vccd1 vccd1 _5441_/X sky130_fd_sc_hd__and2b_1
X_8160_ _8073_/A _8160_/B vssd1 vssd1 vccd1 vccd1 _8160_/X sky130_fd_sc_hd__and2b_1
X_5372_ _8467_/Q _8509_/Q vssd1 vssd1 vccd1 vccd1 _5373_/A sky130_fd_sc_hd__or2b_1
X_4323_ _4326_/A vssd1 vssd1 vccd1 vccd1 _4323_/Y sky130_fd_sc_hd__inv_2
X_7111_ _7153_/A _7111_/B vssd1 vssd1 vccd1 vccd1 _7156_/B sky130_fd_sc_hd__xnor2_1
X_8091_ _8091_/A _8091_/B vssd1 vssd1 vccd1 vccd1 _8111_/A sky130_fd_sc_hd__nand2_1
X_7042_ _7033_/X _7036_/X _7152_/B vssd1 vssd1 vccd1 vccd1 _7099_/B sky130_fd_sc_hd__a21bo_1
XFILLER_67_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7944_ _7944_/A _7944_/B vssd1 vssd1 vccd1 vccd1 _7944_/Y sky130_fd_sc_hd__nand2_1
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7875_ _7868_/A _7875_/B vssd1 vssd1 vccd1 vccd1 _7875_/X sky130_fd_sc_hd__and2b_1
X_6826_ _6826_/A _6870_/A _6826_/C vssd1 vssd1 vccd1 vccd1 _6827_/B sky130_fd_sc_hd__nand3_1
XFILLER_23_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6757_ _6816_/B _6758_/C _6758_/A vssd1 vssd1 vccd1 vccd1 _6879_/C sky130_fd_sc_hd__a21o_1
XFILLER_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5708_ _6244_/B _5689_/A _5706_/A vssd1 vssd1 vccd1 vccd1 _5708_/X sky130_fd_sc_hd__a21o_1
X_6688_ _6688_/A _6781_/B vssd1 vssd1 vccd1 vccd1 _7294_/B sky130_fd_sc_hd__xnor2_2
X_5639_ _5639_/A _5718_/B _5639_/C vssd1 vssd1 vccd1 vccd1 _5669_/A sky130_fd_sc_hd__nand3_1
X_8427_ _8423_/A _7448_/X _8426_/Y _6462_/X vssd1 vssd1 vccd1 vccd1 _8586_/D sky130_fd_sc_hd__a211o_1
X_8358_ _8358_/A _8358_/B vssd1 vssd1 vccd1 vccd1 _8358_/Y sky130_fd_sc_hd__xnor2_1
X_7309_ _7309_/A _7309_/B vssd1 vssd1 vccd1 vccd1 _7313_/A sky130_fd_sc_hd__xnor2_1
XFILLER_2_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8289_ _8346_/A _8289_/B vssd1 vssd1 vccd1 vccd1 _8290_/B sky130_fd_sc_hd__xnor2_1
XFILLER_77_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5990_ _5990_/A _5990_/B _5990_/C vssd1 vssd1 vccd1 vccd1 _5991_/B sky130_fd_sc_hd__nand3_1
XFILLER_91_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4941_ _4987_/A _5071_/A _5164_/A _4941_/D vssd1 vssd1 vccd1 vccd1 _4941_/X sky130_fd_sc_hd__or4_1
XFILLER_17_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4872_ _5053_/B _5138_/B vssd1 vssd1 vccd1 vccd1 _5136_/C sky130_fd_sc_hd__or2_2
XFILLER_17_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7660_ _7660_/A _7660_/B vssd1 vssd1 vccd1 vccd1 _7661_/B sky130_fd_sc_hd__xor2_1
X_6611_ _6640_/B vssd1 vssd1 vccd1 vccd1 _6622_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_7591_ _7888_/A _7742_/A vssd1 vssd1 vccd1 vccd1 _8054_/A sky130_fd_sc_hd__or2_1
XFILLER_32_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6542_ _6609_/B vssd1 vssd1 vccd1 vccd1 _6627_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6473_ _8457_/Q _8561_/Q vssd1 vssd1 vccd1 vccd1 _6486_/A sky130_fd_sc_hd__or2b_1
X_5424_ _6244_/A _5684_/A vssd1 vssd1 vccd1 vccd1 _5522_/A sky130_fd_sc_hd__nand2_1
X_8212_ _8356_/A _8356_/B vssd1 vssd1 vccd1 vccd1 _8212_/X sky130_fd_sc_hd__or2b_1
X_8143_ _8247_/A _8247_/B vssd1 vssd1 vccd1 vccd1 _8248_/B sky130_fd_sc_hd__xor2_1
X_5355_ _5354_/X _5349_/B _5347_/B vssd1 vssd1 vccd1 vccd1 _5357_/C sky130_fd_sc_hd__a21oi_1
X_4306_ _4308_/A vssd1 vssd1 vccd1 vccd1 _4306_/Y sky130_fd_sc_hd__inv_2
XINSDIODE2_6 _7253_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5286_ _8503_/Q _5286_/B vssd1 vssd1 vccd1 vccd1 _5290_/B sky130_fd_sc_hd__and2_1
X_8074_ _8074_/A _8074_/B vssd1 vssd1 vccd1 vccd1 _8133_/B sky130_fd_sc_hd__xor2_1
X_7025_ _7021_/Y _7023_/Y _7024_/X _6961_/B vssd1 vssd1 vccd1 vccd1 _7272_/B sky130_fd_sc_hd__o211ai_2
XFILLER_55_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7927_ _7926_/A _8097_/A _7926_/D _7926_/C vssd1 vssd1 vccd1 vccd1 _7927_/X sky130_fd_sc_hd__a31o_1
XFILLER_36_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7858_ _7618_/A _7615_/B _7618_/C _7613_/X _7583_/A vssd1 vssd1 vccd1 vccd1 _8064_/A
+ sky130_fd_sc_hd__a311o_4
XFILLER_23_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6809_ _6858_/A _6832_/C _6810_/A vssd1 vssd1 vccd1 vccd1 _7296_/A sky130_fd_sc_hd__a21oi_1
XFILLER_23_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7789_ _7788_/A _7788_/B _7788_/C vssd1 vssd1 vccd1 vccd1 _7789_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_23_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8663__79 vssd1 vssd1 vccd1 vccd1 _8663__79/HI _8772_/A sky130_fd_sc_hd__conb_1
XFILLER_65_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5140_ _5174_/S _5109_/B _5134_/X _5139_/X _4623_/X vssd1 vssd1 vccd1 vccd1 _5140_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_69_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5071_ _5071_/A _5099_/C _5071_/C vssd1 vssd1 vccd1 vccd1 _5093_/D sky130_fd_sc_hd__or3_1
XFILLER_69_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8761_ _8761_/A _4344_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[8] sky130_fd_sc_hd__ebufn_8
X_5973_ _5900_/A _5900_/B _5905_/B _5972_/Y vssd1 vssd1 vccd1 vccd1 _6115_/B sky130_fd_sc_hd__a31o_1
XFILLER_37_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4924_ _5164_/A _4920_/X _4921_/X _4977_/C vssd1 vssd1 vccd1 vccd1 _4924_/X sky130_fd_sc_hd__o22a_1
XFILLER_52_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7712_ _8367_/A _7925_/B _7712_/C vssd1 vssd1 vccd1 vccd1 _7712_/X sky130_fd_sc_hd__and3_1
X_8692_ _8692_/A _4269_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[9] sky130_fd_sc_hd__ebufn_8
XFILLER_33_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4855_ _4855_/A vssd1 vssd1 vccd1 vccd1 _5030_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7643_ _8576_/Q _7644_/B vssd1 vssd1 vccd1 vccd1 _7822_/A sky130_fd_sc_hd__or2_1
X_4786_ _4791_/A _4786_/B vssd1 vssd1 vccd1 vccd1 _4956_/C sky130_fd_sc_hd__nor2_1
X_7574_ _7574_/A _7574_/B vssd1 vssd1 vccd1 vccd1 _7607_/A sky130_fd_sc_hd__xnor2_2
X_6525_ _6513_/X _6570_/B _6570_/C _6512_/A _7069_/A vssd1 vssd1 vccd1 vccd1 _6558_/A
+ sky130_fd_sc_hd__a311o_2
X_6456_ _6432_/A _6466_/A _6453_/X _6455_/X vssd1 vssd1 vccd1 vccd1 _8554_/D sky130_fd_sc_hd__a31o_1
X_6387_ _8546_/Q _6386_/A _8547_/Q vssd1 vssd1 vccd1 vccd1 _6387_/Y sky130_fd_sc_hd__a21oi_1
X_5407_ _5694_/A _5579_/B _5408_/C vssd1 vssd1 vccd1 vccd1 _5538_/A sky130_fd_sc_hd__a21oi_1
X_8126_ _8127_/A _8127_/B vssd1 vssd1 vccd1 vccd1 _8257_/A sky130_fd_sc_hd__nor2_1
X_5338_ _5335_/A _5332_/X _5333_/X _5337_/Y vssd1 vssd1 vccd1 vccd1 _8510_/D sky130_fd_sc_hd__a22o_1
X_8057_ _8057_/A _8057_/B vssd1 vssd1 vccd1 vccd1 _8058_/B sky130_fd_sc_hd__or2_1
X_7008_ _7126_/A _7008_/B vssd1 vssd1 vccd1 vccd1 _7075_/A sky130_fd_sc_hd__nor2_2
X_5269_ _6392_/C _5270_/C _5268_/Y vssd1 vssd1 vccd1 vccd1 _8497_/D sky130_fd_sc_hd__a21oi_1
XFILLER_87_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4640_ _4640_/A _5046_/A vssd1 vssd1 vccd1 vccd1 _4640_/Y sky130_fd_sc_hd__nand2_1
XFILLER_30_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6310_ _6362_/B _8535_/Q _6308_/X _6309_/X vssd1 vssd1 vccd1 vccd1 _6310_/X sky130_fd_sc_hd__a31o_1
X_4571_ _8451_/Q _4570_/B _4536_/X vssd1 vssd1 vccd1 vccd1 _4572_/B sky130_fd_sc_hd__o21ai_1
X_7290_ _6893_/A _6846_/B _6854_/B _7289_/X vssd1 vssd1 vccd1 vccd1 _7302_/A sky130_fd_sc_hd__a31o_1
XFILLER_89_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6241_ _6241_/A _6241_/B vssd1 vssd1 vccd1 vccd1 _6241_/X sky130_fd_sc_hd__xor2_1
X_6172_ _6241_/A _6241_/B _6236_/C _6171_/Y _6169_/B vssd1 vssd1 vccd1 vccd1 _6230_/A
+ sky130_fd_sc_hd__a32o_2
X_5123_ _5049_/A _5110_/X _5118_/X _5059_/A _5122_/X vssd1 vssd1 vccd1 vccd1 _5123_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_84_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5054_ _5080_/C _5054_/B vssd1 vssd1 vccd1 vccd1 _5054_/X sky130_fd_sc_hd__or2_1
XFILLER_84_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8744_ _8744_/A _4332_/Y vssd1 vssd1 vccd1 vccd1 io_out[29] sky130_fd_sc_hd__ebufn_8
XFILLER_80_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5956_ _5956_/A _5995_/B vssd1 vssd1 vccd1 vccd1 _5957_/B sky130_fd_sc_hd__xnor2_2
XFILLER_13_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4907_ _5092_/C _4900_/X _4904_/X _4596_/A _4906_/X vssd1 vssd1 vccd1 vccd1 _4907_/X
+ sky130_fd_sc_hd__o221a_1
X_5887_ _5887_/A _5887_/B vssd1 vssd1 vccd1 vccd1 _5888_/B sky130_fd_sc_hd__or2_1
XFILLER_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4838_ _5064_/D vssd1 vssd1 vccd1 vccd1 _5089_/A sky130_fd_sc_hd__clkbuf_2
X_7626_ _7740_/A vssd1 vssd1 vccd1 vccd1 _8146_/A sky130_fd_sc_hd__clkbuf_2
X_4769_ _4886_/A _5156_/A vssd1 vssd1 vccd1 vccd1 _4929_/A sky130_fd_sc_hd__or2_1
X_7557_ _8457_/Q _8581_/Q vssd1 vssd1 vccd1 vccd1 _7569_/A sky130_fd_sc_hd__or2b_2
X_6508_ _7183_/A _7248_/B _6508_/C vssd1 vssd1 vccd1 vccd1 _6509_/B sky130_fd_sc_hd__and3b_1
X_7488_ _7487_/X _7483_/A _7488_/S vssd1 vssd1 vccd1 vccd1 _7489_/B sky130_fd_sc_hd__mux2_1
X_6439_ _6439_/A _6445_/B vssd1 vssd1 vccd1 vccd1 _6440_/B sky130_fd_sc_hd__and2_1
X_8109_ _8238_/B _8109_/B vssd1 vssd1 vccd1 vccd1 _8111_/C sky130_fd_sc_hd__xor2_1
XFILLER_29_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8633__49 vssd1 vssd1 vccd1 vccd1 _8633__49/HI _8742_/A sky130_fd_sc_hd__conb_1
XFILLER_90_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6790_ _6791_/A _6791_/B _6789_/Y vssd1 vssd1 vccd1 vccd1 _6792_/B sky130_fd_sc_hd__o21bai_1
X_5810_ _5870_/A _5810_/B vssd1 vssd1 vccd1 vccd1 _5813_/A sky130_fd_sc_hd__nand2_1
X_5741_ _5785_/A _5785_/B vssd1 vssd1 vccd1 vccd1 _5754_/B sky130_fd_sc_hd__xnor2_1
X_8460_ input3/X _8460_/D vssd1 vssd1 vccd1 vccd1 _8460_/Q sky130_fd_sc_hd__dfxtp_1
X_7411_ _7410_/B _7410_/C _7410_/A vssd1 vssd1 vccd1 vccd1 _7412_/C sky130_fd_sc_hd__o21ai_1
X_5672_ _5669_/X _5670_/Y _5521_/A _5555_/B vssd1 vssd1 vccd1 vccd1 _5673_/C sky130_fd_sc_hd__o211a_1
X_4623_ _5069_/A vssd1 vssd1 vccd1 vccd1 _4623_/X sky130_fd_sc_hd__clkbuf_2
X_8391_ _8391_/A _8568_/Q vssd1 vssd1 vccd1 vccd1 _8392_/B sky130_fd_sc_hd__or2b_1
X_7342_ _7342_/A _7342_/B vssd1 vssd1 vccd1 vccd1 _7342_/Y sky130_fd_sc_hd__xnor2_1
X_4554_ _4557_/C _4554_/B vssd1 vssd1 vccd1 vccd1 _8445_/D sky130_fd_sc_hd__nor2_1
X_7273_ _7097_/B _7271_/X _7272_/X vssd1 vssd1 vccd1 vccd1 _7273_/Y sky130_fd_sc_hd__a21oi_1
X_4485_ _8484_/Q _4491_/B vssd1 vssd1 vccd1 vccd1 _4486_/A sky130_fd_sc_hd__and2_1
XFILLER_89_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6224_ _6224_/A _6165_/B vssd1 vssd1 vccd1 vccd1 _6225_/B sky130_fd_sc_hd__or2b_1
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6155_ _6155_/A _6155_/B vssd1 vssd1 vccd1 vccd1 _6156_/B sky130_fd_sc_hd__or2_1
X_5106_ _5121_/B _4883_/B _5054_/B _5099_/X _5105_/X vssd1 vssd1 vccd1 vccd1 _5107_/D
+ sky130_fd_sc_hd__o221a_1
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6086_ _6086_/A _6086_/B vssd1 vssd1 vccd1 vccd1 _6238_/B sky130_fd_sc_hd__xnor2_2
X_5037_ _5148_/A _5104_/B _4906_/B _5110_/A _4955_/A vssd1 vssd1 vccd1 vccd1 _5037_/X
+ sky130_fd_sc_hd__o41a_1
XFILLER_85_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6988_ _7058_/A _7131_/A vssd1 vssd1 vccd1 vccd1 _6993_/A sky130_fd_sc_hd__nand2_1
X_8727_ _8727_/A _4312_/Y vssd1 vssd1 vccd1 vccd1 io_out[12] sky130_fd_sc_hd__ebufn_8
X_5939_ _6137_/C _5724_/Y _5841_/A _5841_/B vssd1 vssd1 vccd1 vccd1 _5945_/A sky130_fd_sc_hd__a22o_1
XFILLER_40_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7609_ _7744_/A _7609_/B vssd1 vssd1 vccd1 vccd1 _7720_/B sky130_fd_sc_hd__xor2_1
XFILLER_76_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4270_ _4270_/A vssd1 vssd1 vccd1 vccd1 _4270_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7960_ _8317_/A _8326_/A vssd1 vssd1 vccd1 vccd1 _8050_/A sky130_fd_sc_hd__or2_1
XFILLER_82_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6911_ _7280_/B _6911_/B vssd1 vssd1 vccd1 vccd1 _6912_/B sky130_fd_sc_hd__xnor2_1
X_7891_ _7898_/A _7898_/B _7944_/B vssd1 vssd1 vccd1 vccd1 _7945_/C sky130_fd_sc_hd__a21oi_1
XFILLER_35_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6842_ _7043_/A _6842_/B vssd1 vssd1 vccd1 vccd1 _6971_/A sky130_fd_sc_hd__nor2_1
XFILLER_23_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6773_ _6773_/A _6774_/A vssd1 vssd1 vccd1 vccd1 _6886_/B sky130_fd_sc_hd__xor2_1
XFILLER_50_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8512_ input3/X _8512_/D vssd1 vssd1 vccd1 vccd1 _8512_/Q sky130_fd_sc_hd__dfxtp_1
X_5724_ _5724_/A _5825_/B _5825_/C vssd1 vssd1 vccd1 vccd1 _5724_/Y sky130_fd_sc_hd__nor3_1
X_8443_ input3/X _8443_/D vssd1 vssd1 vccd1 vccd1 _8443_/Q sky130_fd_sc_hd__dfxtp_1
X_5655_ _5683_/A _5683_/B vssd1 vssd1 vccd1 vccd1 _5699_/B sky130_fd_sc_hd__xnor2_1
X_4606_ _5162_/A vssd1 vssd1 vccd1 vccd1 _5102_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_8374_ _8369_/X _8373_/X _6261_/X _8577_/Q vssd1 vssd1 vccd1 vccd1 _8577_/D sky130_fd_sc_hd__o2bb2a_1
X_7325_ _6840_/B _7325_/B vssd1 vssd1 vccd1 vccd1 _7325_/X sky130_fd_sc_hd__and2b_1
XFILLER_7_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5586_ _5586_/A _5586_/B vssd1 vssd1 vccd1 vccd1 _6247_/B sky130_fd_sc_hd__xor2_1
XFILLER_89_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4537_ _8440_/Q _4539_/C _4536_/X vssd1 vssd1 vccd1 vccd1 _4537_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_89_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7256_ _7256_/A _7256_/B vssd1 vssd1 vccd1 vccd1 _7256_/Y sky130_fd_sc_hd__nor2_1
X_4468_ _4655_/A _6514_/A vssd1 vssd1 vccd1 vccd1 _4659_/A sky130_fd_sc_hd__nand2_1
X_7187_ _7187_/A _7187_/B _7187_/C vssd1 vssd1 vccd1 vccd1 _7211_/A sky130_fd_sc_hd__and3_1
XFILLER_77_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6207_ _6207_/A _6207_/B vssd1 vssd1 vccd1 vccd1 _6208_/B sky130_fd_sc_hd__nor2_1
X_4399_ _8461_/Q vssd1 vssd1 vccd1 vccd1 _6521_/B sky130_fd_sc_hd__clkbuf_4
X_6138_ _5487_/X _5942_/B _6137_/X vssd1 vssd1 vccd1 vccd1 _6140_/A sky130_fd_sc_hd__o21a_1
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8603__19 vssd1 vssd1 vccd1 vccd1 _8603__19/HI _8698_/A sky130_fd_sc_hd__conb_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6069_ _6079_/A _6069_/B vssd1 vssd1 vccd1 vccd1 _6069_/X sky130_fd_sc_hd__xor2_1
XFILLER_73_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5440_ _8521_/Q _7559_/B vssd1 vssd1 vccd1 vccd1 _5455_/B sky130_fd_sc_hd__xnor2_2
X_5371_ _5371_/A vssd1 vssd1 vccd1 vccd1 _8515_/D sky130_fd_sc_hd__clkbuf_1
X_8669__85 vssd1 vssd1 vccd1 vccd1 _8669__85/HI _8778_/A sky130_fd_sc_hd__conb_1
X_4322_ _4326_/A vssd1 vssd1 vccd1 vccd1 _4322_/Y sky130_fd_sc_hd__inv_2
X_7110_ _7129_/A _7129_/B vssd1 vssd1 vccd1 vccd1 _7111_/B sky130_fd_sc_hd__xnor2_1
X_8090_ _8046_/A _8046_/B _8047_/B _8047_/A vssd1 vssd1 vccd1 vccd1 _8114_/A sky130_fd_sc_hd__o2bb2ai_4
X_7041_ _7101_/A _7102_/A _7040_/Y vssd1 vssd1 vccd1 vccd1 _7152_/B sky130_fd_sc_hd__o21ai_2
XFILLER_79_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7943_ _7903_/A _7903_/B _7942_/Y vssd1 vssd1 vccd1 vccd1 _8048_/A sky130_fd_sc_hd__o21ai_2
X_7874_ _8180_/A _8180_/B _7873_/X vssd1 vssd1 vccd1 vccd1 _7937_/B sky130_fd_sc_hd__a21o_1
X_6825_ _6826_/A _6870_/A _6826_/C vssd1 vssd1 vccd1 vccd1 _6825_/Y sky130_fd_sc_hd__a21oi_1
X_6756_ _6875_/B _6875_/A vssd1 vssd1 vccd1 vccd1 _6758_/A sky130_fd_sc_hd__and2b_1
XFILLER_50_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5707_ _5581_/A _6183_/S _5992_/A vssd1 vssd1 vccd1 vccd1 _5707_/Y sky130_fd_sc_hd__o21ai_1
X_6687_ _6687_/A vssd1 vssd1 vccd1 vccd1 _6781_/B sky130_fd_sc_hd__buf_2
XFILLER_12_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8426_ _8426_/A _8426_/B vssd1 vssd1 vccd1 vccd1 _8426_/Y sky130_fd_sc_hd__nor2_1
X_5638_ _5637_/A _5637_/B _5718_/A _5636_/X vssd1 vssd1 vccd1 vccd1 _5639_/C sky130_fd_sc_hd__a2bb2o_1
X_8357_ _8361_/A _8361_/B _8213_/X vssd1 vssd1 vccd1 vccd1 _8358_/B sky130_fd_sc_hd__a21o_1
X_5569_ _5738_/A vssd1 vssd1 vccd1 vccd1 _5839_/A sky130_fd_sc_hd__clkbuf_2
X_7308_ _7308_/A _7308_/B vssd1 vssd1 vccd1 vccd1 _7309_/B sky130_fd_sc_hd__xnor2_1
XFILLER_2_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8288_ _8288_/A _8345_/A vssd1 vssd1 vccd1 vccd1 _8289_/B sky130_fd_sc_hd__xnor2_1
X_7239_ _7239_/A _7253_/A vssd1 vssd1 vccd1 vccd1 _7240_/A sky130_fd_sc_hd__nor2_1
XFILLER_77_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4940_ _5153_/A _5112_/B vssd1 vssd1 vccd1 vccd1 _4941_/D sky130_fd_sc_hd__or2_1
XFILLER_45_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4871_ _4871_/A vssd1 vssd1 vccd1 vccd1 _5053_/B sky130_fd_sc_hd__clkbuf_2
X_6610_ _6627_/B _6627_/C _6627_/A vssd1 vssd1 vccd1 vccd1 _6640_/B sky130_fd_sc_hd__a21oi_1
X_7590_ _7607_/A vssd1 vssd1 vccd1 vccd1 _7742_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_32_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6541_ _6541_/A _7539_/B vssd1 vssd1 vccd1 vccd1 _6609_/B sky130_fd_sc_hd__nand2_1
XFILLER_9_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6472_ _7412_/A vssd1 vssd1 vccd1 vccd1 _6472_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_9_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5423_ _5532_/A _5532_/B vssd1 vssd1 vccd1 vccd1 _5684_/A sky130_fd_sc_hd__xor2_4
X_8211_ _8211_/A _8211_/B vssd1 vssd1 vccd1 vccd1 _8356_/B sky130_fd_sc_hd__xor2_1
X_5354_ _5360_/B _5345_/B vssd1 vssd1 vccd1 vccd1 _5354_/X sky130_fd_sc_hd__or2b_1
X_8142_ _8142_/A _8142_/B vssd1 vssd1 vccd1 vccd1 _8247_/B sky130_fd_sc_hd__xnor2_1
X_4305_ _4308_/A vssd1 vssd1 vccd1 vccd1 _4305_/Y sky130_fd_sc_hd__inv_2
XFILLER_87_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_7 _7253_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5285_ _5286_/B _5285_/B vssd1 vssd1 vccd1 vccd1 _8502_/D sky130_fd_sc_hd__nor2_1
X_8073_ _8073_/A _8160_/B vssd1 vssd1 vccd1 vccd1 _8074_/B sky130_fd_sc_hd__xnor2_1
X_7024_ _6961_/A _6960_/C _6960_/B vssd1 vssd1 vccd1 vccd1 _7024_/X sky130_fd_sc_hd__a21o_1
XFILLER_59_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7926_ _7926_/A _8097_/A _7926_/C _7926_/D vssd1 vssd1 vccd1 vccd1 _8003_/A sky130_fd_sc_hd__and4_1
XFILLER_70_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7857_ _7877_/B _7878_/B vssd1 vssd1 vccd1 vccd1 _7867_/A sky130_fd_sc_hd__xnor2_1
X_6808_ _7032_/B _7032_/C _6806_/A vssd1 vssd1 vccd1 vccd1 _6832_/C sky130_fd_sc_hd__a21oi_2
XFILLER_23_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7788_ _7788_/A _7788_/B _7788_/C vssd1 vssd1 vccd1 vccd1 _7788_/X sky130_fd_sc_hd__and3_1
X_6739_ _6739_/A _6739_/B _6736_/X vssd1 vssd1 vccd1 vccd1 _6802_/C sky130_fd_sc_hd__or3b_2
X_8409_ _8408_/Y _8405_/A _8430_/A vssd1 vssd1 vccd1 vccd1 _8410_/B sky130_fd_sc_hd__mux2_1
XFILLER_78_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8639__55 vssd1 vssd1 vccd1 vccd1 _8639__55/HI _8748_/A sky130_fd_sc_hd__conb_1
XFILLER_89_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5070_ _4808_/A _4817_/A _4953_/B vssd1 vssd1 vccd1 vccd1 _5173_/A sky130_fd_sc_hd__a21oi_2
XFILLER_84_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8760_ _8760_/A _4342_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[7] sky130_fd_sc_hd__ebufn_8
XFILLER_52_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5972_ _6226_/A _5972_/B vssd1 vssd1 vccd1 vccd1 _5972_/Y sky130_fd_sc_hd__nor2_1
X_4923_ _5093_/A _5087_/B vssd1 vssd1 vccd1 vccd1 _4977_/C sky130_fd_sc_hd__or2_1
XFILLER_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7711_ _7822_/B vssd1 vssd1 vccd1 vccd1 _7925_/B sky130_fd_sc_hd__clkbuf_2
X_8691_ _8691_/A _4268_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[8] sky130_fd_sc_hd__ebufn_8
XFILLER_33_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4854_ _5036_/A _5093_/B vssd1 vssd1 vccd1 vccd1 _5148_/B sky130_fd_sc_hd__or2_1
XFILLER_20_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7642_ _8099_/A _7978_/A vssd1 vssd1 vccd1 vccd1 _7658_/B sky130_fd_sc_hd__nor2_1
X_4785_ _4792_/A _4786_/B vssd1 vssd1 vccd1 vccd1 _5162_/B sky130_fd_sc_hd__nor2_2
XFILLER_20_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7573_ _8052_/A vssd1 vssd1 vccd1 vccd1 _7756_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6524_ _6524_/A vssd1 vssd1 vccd1 vccd1 _6570_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_6455_ _6455_/A _7399_/B _7406_/A vssd1 vssd1 vccd1 vccd1 _6455_/X sky130_fd_sc_hd__and3_1
X_6386_ _6386_/A _6386_/B vssd1 vssd1 vccd1 vccd1 _8545_/D sky130_fd_sc_hd__nor2_1
X_5406_ _5651_/A _5406_/B vssd1 vssd1 vccd1 vccd1 _5408_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8125_ _8125_/A _8125_/B vssd1 vssd1 vccd1 vccd1 _8127_/B sky130_fd_sc_hd__xnor2_1
X_5337_ _8509_/Q _5337_/B vssd1 vssd1 vccd1 vccd1 _5337_/Y sky130_fd_sc_hd__xnor2_1
X_5268_ _6392_/C _5270_/C _5230_/B vssd1 vssd1 vccd1 vccd1 _5268_/Y sky130_fd_sc_hd__o21ai_1
X_8056_ _8057_/A _8057_/B vssd1 vssd1 vccd1 vccd1 _8129_/A sky130_fd_sc_hd__nand2_1
X_7007_ _7007_/A _7055_/A vssd1 vssd1 vccd1 vccd1 _7008_/B sky130_fd_sc_hd__xnor2_1
X_5199_ _8478_/Q _5205_/B vssd1 vssd1 vccd1 vccd1 _5199_/X sky130_fd_sc_hd__or2_1
XFILLER_75_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7909_ _7909_/A _7909_/B vssd1 vssd1 vccd1 vccd1 _7939_/B sky130_fd_sc_hd__xor2_2
XFILLER_70_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4570_ _8451_/Q _4570_/B vssd1 vssd1 vccd1 vccd1 _4574_/B sky130_fd_sc_hd__and2_1
XFILLER_6_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6240_ _6069_/X _6231_/Y _6232_/Y _6235_/Y _6239_/X vssd1 vssd1 vccd1 vccd1 _6240_/Y
+ sky130_fd_sc_hd__o2111ai_1
XFILLER_6_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6171_ _6236_/A _6236_/B _6169_/A vssd1 vssd1 vccd1 vccd1 _6171_/Y sky130_fd_sc_hd__o21ai_1
X_5122_ _4955_/A _5116_/B _5002_/D _5117_/X vssd1 vssd1 vccd1 vccd1 _5122_/X sky130_fd_sc_hd__a211o_1
XFILLER_69_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5053_ _5162_/A _5053_/B vssd1 vssd1 vccd1 vccd1 _5054_/B sky130_fd_sc_hd__or2_1
XFILLER_65_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8743_ _8743_/A _4331_/Y vssd1 vssd1 vccd1 vccd1 io_out[28] sky130_fd_sc_hd__ebufn_8
XFILLER_80_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5955_ _5955_/A _6013_/B vssd1 vssd1 vccd1 vccd1 _5995_/B sky130_fd_sc_hd__xnor2_2
XFILLER_40_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4906_ _4956_/C _4906_/B _5059_/A _4906_/D vssd1 vssd1 vccd1 vccd1 _4906_/X sky130_fd_sc_hd__or4_1
XFILLER_52_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5886_ _5887_/A _5887_/B vssd1 vssd1 vccd1 vccd1 _5888_/A sky130_fd_sc_hd__nand2_1
X_4837_ _4973_/A vssd1 vssd1 vccd1 vccd1 _4839_/A sky130_fd_sc_hd__clkbuf_2
X_7625_ _7725_/C vssd1 vssd1 vccd1 vccd1 _8147_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_21_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4768_ _4706_/C _4756_/A _4943_/B _4767_/Y vssd1 vssd1 vccd1 vccd1 _5156_/A sky130_fd_sc_hd__a211o_2
X_7556_ _7556_/A _7556_/B vssd1 vssd1 vccd1 vccd1 _7574_/A sky130_fd_sc_hd__nor2_2
X_6507_ _6507_/A vssd1 vssd1 vccd1 vccd1 _7248_/B sky130_fd_sc_hd__clkbuf_2
X_4699_ _5370_/A _4699_/B _4702_/B vssd1 vssd1 vccd1 vccd1 _4700_/A sky130_fd_sc_hd__and3_1
X_7487_ _8574_/Q _7487_/B vssd1 vssd1 vccd1 vccd1 _7487_/X sky130_fd_sc_hd__or2_1
XFILLER_20_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6438_ _6439_/A _6445_/B vssd1 vssd1 vccd1 vccd1 _6440_/A sky130_fd_sc_hd__nor2_1
X_6369_ _6371_/B _6371_/C _6331_/B vssd1 vssd1 vccd1 vccd1 _6369_/Y sky130_fd_sc_hd__o21ai_1
X_8108_ _8108_/A _8108_/B vssd1 vssd1 vccd1 vccd1 _8109_/B sky130_fd_sc_hd__xnor2_1
XFILLER_29_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8039_ _8039_/A _7977_/B vssd1 vssd1 vccd1 vccd1 _8039_/X sky130_fd_sc_hd__or2b_1
XFILLER_75_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8609__25 vssd1 vssd1 vccd1 vccd1 _8609__25/HI _8704_/A sky130_fd_sc_hd__conb_1
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5740_ _5824_/A _5740_/B vssd1 vssd1 vccd1 vccd1 _5785_/B sky130_fd_sc_hd__xnor2_1
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7410_ _7410_/A _7410_/B _7410_/C vssd1 vssd1 vccd1 vccd1 _7412_/B sky130_fd_sc_hd__or3_1
X_5671_ _5521_/A _5555_/B _5669_/X _5670_/Y vssd1 vssd1 vccd1 vccd1 _5673_/B sky130_fd_sc_hd__a211oi_1
X_4622_ _4629_/A _4621_/Y _4657_/B vssd1 vssd1 vccd1 vccd1 _8456_/D sky130_fd_sc_hd__a21boi_1
XFILLER_30_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8390_ _8568_/Q _8391_/A vssd1 vssd1 vccd1 vccd1 _8392_/A sky130_fd_sc_hd__or2b_1
X_7341_ _7258_/Y _7341_/B vssd1 vssd1 vccd1 vccd1 _7342_/B sky130_fd_sc_hd__and2b_1
X_4553_ _8445_/Q _4552_/B _4536_/X vssd1 vssd1 vccd1 vccd1 _4554_/B sky130_fd_sc_hd__o21ai_1
X_4484_ _4484_/A vssd1 vssd1 vccd1 vccd1 _8737_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7272_ _7272_/A _7272_/B _7272_/C vssd1 vssd1 vccd1 vccd1 _7272_/X sky130_fd_sc_hd__and3_1
XFILLER_89_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6223_ _6223_/A _6164_/B vssd1 vssd1 vccd1 vccd1 _6225_/A sky130_fd_sc_hd__or2b_1
XFILLER_85_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6154_ _6154_/A _6154_/B vssd1 vssd1 vccd1 vccd1 _6155_/B sky130_fd_sc_hd__and2_1
X_5105_ _4977_/C _5104_/X _8455_/Q _5030_/B vssd1 vssd1 vccd1 vccd1 _5105_/X sky130_fd_sc_hd__a211o_1
XFILLER_85_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6085_ _6087_/A _6090_/C vssd1 vssd1 vccd1 vccd1 _6086_/B sky130_fd_sc_hd__xor2_1
X_5036_ _5036_/A _5147_/B vssd1 vssd1 vccd1 vccd1 _5110_/A sky130_fd_sc_hd__or2_1
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6987_ _7118_/A _6987_/B vssd1 vssd1 vccd1 vccd1 _7131_/A sky130_fd_sc_hd__xnor2_4
X_8726_ _8726_/A _4311_/Y vssd1 vssd1 vccd1 vccd1 io_out[11] sky130_fd_sc_hd__ebufn_8
XFILLER_15_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5938_ _5938_/A _6025_/B vssd1 vssd1 vccd1 vccd1 _6137_/C sky130_fd_sc_hd__nor2_2
XFILLER_80_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5869_ _5870_/A _5870_/B vssd1 vssd1 vccd1 vccd1 _5871_/A sky130_fd_sc_hd__or2_1
X_7608_ _7607_/Y _7607_/B _7725_/A vssd1 vssd1 vccd1 vccd1 _7609_/B sky130_fd_sc_hd__mux2_1
X_7539_ _7539_/A _7539_/B vssd1 vssd1 vccd1 vccd1 _7539_/Y sky130_fd_sc_hd__nand2_1
XFILLER_48_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6910_ _6909_/A _6910_/B vssd1 vssd1 vccd1 vccd1 _6911_/B sky130_fd_sc_hd__and2b_1
X_7890_ _7898_/A _7898_/B _7944_/B vssd1 vssd1 vccd1 vccd1 _7945_/B sky130_fd_sc_hd__and3_1
X_6841_ _6837_/A _6836_/C _6836_/A vssd1 vssd1 vccd1 vccd1 _6848_/B sky130_fd_sc_hd__a21o_1
XFILLER_22_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6772_ _6828_/A _6772_/B vssd1 vssd1 vccd1 vccd1 _6774_/A sky130_fd_sc_hd__or2_1
X_8511_ input3/X _8511_/D vssd1 vssd1 vccd1 vccd1 _8511_/Q sky130_fd_sc_hd__dfxtp_1
X_5723_ _5767_/A _5767_/B vssd1 vssd1 vccd1 vccd1 _5765_/A sky130_fd_sc_hd__nor2_2
X_5654_ _5659_/A _5685_/C vssd1 vssd1 vccd1 vccd1 _5683_/B sky130_fd_sc_hd__xnor2_1
XFILLER_30_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8442_ input3/X _8442_/D vssd1 vssd1 vccd1 vccd1 _8442_/Q sky130_fd_sc_hd__dfxtp_1
X_4605_ _5001_/A vssd1 vssd1 vccd1 vccd1 _5162_/A sky130_fd_sc_hd__clkbuf_2
X_8373_ _8385_/B _8385_/C _8372_/Y _7399_/B vssd1 vssd1 vccd1 vccd1 _8373_/X sky130_fd_sc_hd__o31a_1
XFILLER_30_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7324_ _7324_/A _7324_/B vssd1 vssd1 vccd1 vccd1 _7330_/A sky130_fd_sc_hd__xnor2_1
X_5585_ _6243_/A _6243_/B vssd1 vssd1 vccd1 vccd1 _6247_/A sky130_fd_sc_hd__or2_1
X_4536_ _4536_/A vssd1 vssd1 vccd1 vccd1 _4536_/X sky130_fd_sc_hd__clkbuf_2
X_7255_ _7349_/A _7349_/B _7243_/A vssd1 vssd1 vccd1 vccd1 _7354_/B sky130_fd_sc_hd__a21o_1
X_4467_ _5526_/B _4706_/A _4467_/C _4591_/C vssd1 vssd1 vccd1 vccd1 _4469_/B sky130_fd_sc_hd__or4_1
X_7186_ _7186_/A _7186_/B vssd1 vssd1 vccd1 vccd1 _7187_/C sky130_fd_sc_hd__xnor2_1
X_4398_ _7575_/B _4638_/A vssd1 vssd1 vccd1 vccd1 _4593_/A sky130_fd_sc_hd__or2_1
X_6206_ _5940_/A _5930_/B _6152_/A _6205_/X vssd1 vssd1 vccd1 vccd1 _6207_/B sky130_fd_sc_hd__o31a_1
X_6137_ _6137_/A _6137_/B _6137_/C vssd1 vssd1 vccd1 vccd1 _6137_/X sky130_fd_sc_hd__or3_1
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6068_ _6170_/A _6068_/B vssd1 vssd1 vccd1 vccd1 _6069_/B sky130_fd_sc_hd__nor2_1
X_5019_ _5019_/A _5019_/B _5104_/C vssd1 vssd1 vccd1 vccd1 _5020_/D sky130_fd_sc_hd__or3_1
XFILLER_26_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8709_ _8709_/A _4291_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[26] sky130_fd_sc_hd__ebufn_8
XFILLER_13_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5370_ _5370_/A _5370_/B _5370_/C vssd1 vssd1 vccd1 vccd1 _5371_/A sky130_fd_sc_hd__and3_1
X_4321_ _4327_/A vssd1 vssd1 vccd1 vccd1 _4326_/A sky130_fd_sc_hd__clkbuf_2
X_7040_ _7038_/A _7038_/B _7180_/B vssd1 vssd1 vccd1 vccd1 _7040_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_67_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7942_ _7942_/A _7942_/B vssd1 vssd1 vccd1 vccd1 _7942_/Y sky130_fd_sc_hd__nand2_1
XFILLER_82_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7873_ _7870_/B _7873_/B vssd1 vssd1 vccd1 vccd1 _7873_/X sky130_fd_sc_hd__and2b_1
X_6824_ _6824_/A _6824_/B vssd1 vssd1 vccd1 vccd1 _6826_/C sky130_fd_sc_hd__xnor2_2
XFILLER_63_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6755_ _6755_/A _6755_/B vssd1 vssd1 vccd1 vccd1 _6875_/A sky130_fd_sc_hd__nand2_1
XFILLER_11_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5706_ _5706_/A vssd1 vssd1 vccd1 vccd1 _5992_/A sky130_fd_sc_hd__buf_2
X_6686_ _6680_/A _7005_/B _6686_/C vssd1 vssd1 vccd1 vccd1 _6687_/A sky130_fd_sc_hd__and3b_1
XFILLER_12_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8425_ _8425_/A _8425_/B vssd1 vssd1 vccd1 vccd1 _8426_/B sky130_fd_sc_hd__xnor2_1
XFILLER_12_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5637_ _5637_/A _5637_/B _5718_/A _5636_/X vssd1 vssd1 vccd1 vccd1 _5718_/B sky130_fd_sc_hd__or4bb_1
X_8356_ _8356_/A _8356_/B vssd1 vssd1 vccd1 vccd1 _8358_/A sky130_fd_sc_hd__xnor2_1
X_5568_ _5764_/A vssd1 vssd1 vccd1 vccd1 _5738_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_88_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7307_ _7293_/A _7039_/B _6857_/B _7306_/X vssd1 vssd1 vccd1 vccd1 _7308_/B sky130_fd_sc_hd__o31a_1
X_8287_ _8287_/A _8297_/B vssd1 vssd1 vccd1 vccd1 _8345_/A sky130_fd_sc_hd__xor2_1
X_4519_ _8434_/Q _8433_/Q _8435_/Q vssd1 vssd1 vccd1 vccd1 _4520_/C sky130_fd_sc_hd__a21o_1
X_7238_ _7244_/A _7244_/B vssd1 vssd1 vccd1 vccd1 _7253_/A sky130_fd_sc_hd__and2_1
X_5499_ _5499_/A _5499_/B _5499_/C vssd1 vssd1 vccd1 vccd1 _5764_/B sky130_fd_sc_hd__and3_1
XFILLER_77_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7169_ _7345_/A _7345_/B _7345_/C vssd1 vssd1 vccd1 vccd1 _7171_/A sky130_fd_sc_hd__or3_1
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4870_ _5039_/B vssd1 vssd1 vccd1 vccd1 _4955_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_60_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6540_ _6609_/A vssd1 vssd1 vccd1 vccd1 _6627_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6471_ _6471_/A vssd1 vssd1 vccd1 vccd1 _8556_/D sky130_fd_sc_hd__clkbuf_1
X_8210_ _8210_/A _8213_/C vssd1 vssd1 vccd1 vccd1 _8356_/A sky130_fd_sc_hd__and2_1
X_5422_ _5422_/A _5422_/B vssd1 vssd1 vccd1 vccd1 _5532_/B sky130_fd_sc_hd__and2_2
X_5353_ _8513_/Q _5359_/B vssd1 vssd1 vccd1 vccd1 _5357_/B sky130_fd_sc_hd__or2b_1
X_8141_ _8141_/A _8141_/B vssd1 vssd1 vccd1 vccd1 _8142_/B sky130_fd_sc_hd__nand2_1
X_4304_ _4308_/A vssd1 vssd1 vccd1 vccd1 _4304_/Y sky130_fd_sc_hd__inv_2
X_5284_ _8502_/Q _5282_/A _5264_/X vssd1 vssd1 vccd1 vccd1 _5285_/B sky130_fd_sc_hd__o21ai_1
X_8072_ _8072_/A _8276_/B vssd1 vssd1 vccd1 vccd1 _8160_/B sky130_fd_sc_hd__xnor2_1
X_7023_ _7017_/B _7019_/C _7021_/Y _7022_/X vssd1 vssd1 vccd1 vccd1 _7023_/Y sky130_fd_sc_hd__a211oi_2
XINSDIODE2_8 _7253_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7925_ _7983_/B _7925_/B vssd1 vssd1 vccd1 vccd1 _7926_/D sky130_fd_sc_hd__or2_1
XFILLER_43_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7856_ _7856_/A _7856_/B vssd1 vssd1 vccd1 vccd1 _7878_/B sky130_fd_sc_hd__xnor2_1
X_6807_ _6810_/B vssd1 vssd1 vccd1 vccd1 _6858_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_23_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4999_ _5151_/A _5132_/C _4988_/X _5004_/C _4998_/X vssd1 vssd1 vccd1 vccd1 _5006_/C
+ sky130_fd_sc_hd__o41a_1
X_7787_ _8198_/A _7787_/B vssd1 vssd1 vccd1 vccd1 _7788_/C sky130_fd_sc_hd__nor2_2
X_6738_ _7033_/A _6736_/B _6806_/A vssd1 vssd1 vccd1 vccd1 _6739_/B sky130_fd_sc_hd__a21o_1
XFILLER_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6669_ _6678_/B _6669_/B vssd1 vssd1 vccd1 vccd1 _6703_/B sky130_fd_sc_hd__xnor2_1
X_8408_ _8408_/A _8414_/B vssd1 vssd1 vccd1 vccd1 _8408_/Y sky130_fd_sc_hd__xnor2_1
X_8339_ _8339_/A _8284_/A vssd1 vssd1 vccd1 vccd1 _8339_/X sky130_fd_sc_hd__or2b_1
XFILLER_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5971_ _5971_/A _5908_/B vssd1 vssd1 vccd1 vccd1 _5990_/B sky130_fd_sc_hd__or2b_1
X_4922_ _5020_/C _4996_/A vssd1 vssd1 vccd1 vccd1 _5087_/B sky130_fd_sc_hd__or2_2
X_8690_ _8690_/A _4267_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[7] sky130_fd_sc_hd__ebufn_8
XFILLER_52_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7710_ _7783_/A vssd1 vssd1 vccd1 vccd1 _7710_/Y sky130_fd_sc_hd__inv_2
X_7641_ _7641_/A _7641_/B vssd1 vssd1 vccd1 vccd1 _8099_/A sky130_fd_sc_hd__xnor2_2
X_4853_ _4944_/B _4899_/B vssd1 vssd1 vccd1 vccd1 _5093_/B sky130_fd_sc_hd__nor2_2
X_4784_ _5087_/A vssd1 vssd1 vccd1 vccd1 _5064_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_7572_ _7620_/A vssd1 vssd1 vccd1 vccd1 _8052_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6523_ _6574_/B _6575_/B _6575_/C _6521_/X _6522_/X vssd1 vssd1 vccd1 vccd1 _6524_/A
+ sky130_fd_sc_hd__a311o_1
XFILLER_20_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6454_ _6465_/A vssd1 vssd1 vccd1 vccd1 _7406_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5405_ _5408_/B vssd1 vssd1 vccd1 vccd1 _5579_/B sky130_fd_sc_hd__clkbuf_2
X_6385_ _8545_/Q _6384_/B _6326_/B vssd1 vssd1 vccd1 vccd1 _6386_/B sky130_fd_sc_hd__o21ai_1
X_8124_ _8227_/A _8348_/A vssd1 vssd1 vccd1 vccd1 _8125_/B sky130_fd_sc_hd__xor2_1
X_5336_ _5336_/A _5336_/B vssd1 vssd1 vccd1 vccd1 _5337_/B sky130_fd_sc_hd__nand2_1
XFILLER_87_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5267_ _8497_/Q vssd1 vssd1 vccd1 vccd1 _6392_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_8055_ _8319_/A _8323_/A _8248_/A vssd1 vssd1 vccd1 vccd1 _8057_/B sky130_fd_sc_hd__o21ba_1
X_7006_ _7122_/C _7116_/B _7148_/B _7005_/X vssd1 vssd1 vccd1 vccd1 _7126_/A sky130_fd_sc_hd__o31a_1
X_5198_ _8519_/Q _5188_/X _5197_/X _6426_/A vssd1 vssd1 vccd1 vccd1 _8477_/D sky130_fd_sc_hd__o211a_1
XFILLER_68_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7908_ _8054_/B _7865_/A _7991_/A vssd1 vssd1 vccd1 vccd1 _7909_/B sky130_fd_sc_hd__a21oi_2
XFILLER_43_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7839_ _7752_/A _7839_/B vssd1 vssd1 vccd1 vccd1 _7868_/A sky130_fd_sc_hd__and2b_1
XFILLER_34_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6170_ _6170_/A vssd1 vssd1 vccd1 vccd1 _6236_/A sky130_fd_sc_hd__inv_2
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5121_ _5121_/A _5121_/B vssd1 vssd1 vccd1 vccd1 _5121_/X sky130_fd_sc_hd__or2_1
X_5052_ _5058_/C vssd1 vssd1 vccd1 vccd1 _5080_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_37_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8742_ _8742_/A _4330_/Y vssd1 vssd1 vccd1 vccd1 io_out[27] sky130_fd_sc_hd__ebufn_8
XFILLER_92_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5954_ _5954_/A _6012_/B vssd1 vssd1 vccd1 vccd1 _6013_/B sky130_fd_sc_hd__xnor2_1
X_4905_ _5162_/A _5019_/A vssd1 vssd1 vccd1 vccd1 _5059_/A sky130_fd_sc_hd__nand2_1
X_5885_ _5914_/B _5885_/B vssd1 vssd1 vccd1 vccd1 _5887_/B sky130_fd_sc_hd__xnor2_1
X_4836_ _5019_/A vssd1 vssd1 vccd1 vccd1 _4973_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_21_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7624_ _7718_/A _7624_/B vssd1 vssd1 vccd1 vccd1 _7633_/A sky130_fd_sc_hd__xnor2_1
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7555_ _7554_/B _8583_/Q vssd1 vssd1 vccd1 vccd1 _7556_/B sky130_fd_sc_hd__and2b_1
X_6506_ _6506_/A vssd1 vssd1 vccd1 vccd1 _6507_/A sky130_fd_sc_hd__inv_2
X_4767_ _4767_/A _4817_/A vssd1 vssd1 vccd1 vccd1 _4767_/Y sky130_fd_sc_hd__nor2_1
X_4698_ _4698_/A _4698_/B _4698_/C vssd1 vssd1 vccd1 vccd1 _4702_/B sky130_fd_sc_hd__nand3_1
X_7486_ _7539_/A _7448_/X _7485_/Y _6462_/X vssd1 vssd1 vccd1 vccd1 _8575_/D sky130_fd_sc_hd__a211o_1
XFILLER_20_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6437_ _6433_/A _5294_/X _6432_/X _6436_/X vssd1 vssd1 vccd1 vccd1 _8551_/D sky130_fd_sc_hd__a22o_1
XFILLER_20_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6368_ _6371_/C _6368_/B vssd1 vssd1 vccd1 vccd1 _8539_/D sky130_fd_sc_hd__nor2_1
XFILLER_96_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8107_ _8249_/A _8107_/B vssd1 vssd1 vccd1 vccd1 _8108_/B sky130_fd_sc_hd__xnor2_1
X_5319_ _8508_/Q vssd1 vssd1 vccd1 vccd1 _5360_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6299_ _5326_/B _6298_/X _8526_/Q vssd1 vssd1 vccd1 vccd1 _6301_/A sky130_fd_sc_hd__a21oi_1
X_8038_ _8038_/A _8038_/B vssd1 vssd1 vccd1 vccd1 _8080_/A sky130_fd_sc_hd__xnor2_1
XFILLER_29_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5670_ _5669_/A _5669_/B _5669_/C vssd1 vssd1 vccd1 vccd1 _5670_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4621_ _5179_/A _4640_/A vssd1 vssd1 vccd1 vccd1 _4621_/Y sky130_fd_sc_hd__nand2_1
XFILLER_30_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7340_ _7217_/Y _7344_/B _7343_/A vssd1 vssd1 vccd1 vccd1 _7342_/A sky130_fd_sc_hd__a21o_1
X_4552_ _8445_/Q _4552_/B vssd1 vssd1 vccd1 vccd1 _4557_/C sky130_fd_sc_hd__and2_1
X_4483_ _8483_/Q _4491_/B vssd1 vssd1 vccd1 vccd1 _4484_/A sky130_fd_sc_hd__and2_1
X_7271_ _7272_/A _7030_/B vssd1 vssd1 vccd1 vccd1 _7271_/X sky130_fd_sc_hd__or2b_1
X_6222_ _6222_/A _6222_/B vssd1 vssd1 vccd1 vccd1 _6227_/A sky130_fd_sc_hd__xnor2_1
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6153_ _6154_/A _6153_/B _6153_/C vssd1 vssd1 vccd1 vccd1 _6155_/A sky130_fd_sc_hd__and3b_1
X_5104_ _5104_/A _5104_/B _5104_/C _5104_/D vssd1 vssd1 vccd1 vccd1 _5104_/X sky130_fd_sc_hd__or4_1
XFILLER_85_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6084_ _6084_/A _6084_/B vssd1 vssd1 vccd1 vccd1 _6090_/C sky130_fd_sc_hd__xor2_1
XFILLER_85_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5035_ _5171_/B _5132_/D _5153_/B _5035_/D vssd1 vssd1 vccd1 vccd1 _5091_/A sky130_fd_sc_hd__or4_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6986_ _7233_/B _6643_/D _6971_/B _6913_/A vssd1 vssd1 vccd1 vccd1 _7058_/A sky130_fd_sc_hd__o22ai_4
X_8725_ _8725_/A _4310_/Y vssd1 vssd1 vccd1 vccd1 io_out[10] sky130_fd_sc_hd__ebufn_8
X_5937_ _5835_/X _5844_/B _5836_/A vssd1 vssd1 vccd1 vccd1 _5954_/A sky130_fd_sc_hd__a21oi_1
XFILLER_15_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5868_ _5868_/A _5868_/B vssd1 vssd1 vccd1 vccd1 _5870_/B sky130_fd_sc_hd__xnor2_1
X_7607_ _7607_/A _7607_/B vssd1 vssd1 vccd1 vccd1 _7607_/Y sky130_fd_sc_hd__xnor2_1
X_4819_ _4676_/A _4953_/A _4798_/B vssd1 vssd1 vccd1 vccd1 _4906_/B sky130_fd_sc_hd__a21oi_4
X_5799_ _6108_/A vssd1 vssd1 vccd1 vccd1 _5918_/C sky130_fd_sc_hd__clkbuf_2
X_8587_ input3/X _8587_/D vssd1 vssd1 vccd1 vccd1 _8587_/Q sky130_fd_sc_hd__dfxtp_1
X_7538_ _8575_/Q _7538_/B vssd1 vssd1 vccd1 vccd1 _7540_/A sky130_fd_sc_hd__nor2_2
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7469_ _8418_/S vssd1 vssd1 vccd1 vccd1 _8426_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_76_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6840_ _7325_/B _6840_/B vssd1 vssd1 vccd1 vccd1 _6862_/A sky130_fd_sc_hd__xnor2_2
XFILLER_35_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6771_ _6771_/A _6771_/B vssd1 vssd1 vccd1 vccd1 _6772_/B sky130_fd_sc_hd__and2_1
XFILLER_35_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5722_ _5722_/A _5722_/B vssd1 vssd1 vccd1 vccd1 _5758_/A sky130_fd_sc_hd__nand2_1
X_8510_ input3/X _8510_/D vssd1 vssd1 vccd1 vccd1 _8510_/Q sky130_fd_sc_hd__dfxtp_2
X_5653_ _6053_/A _5653_/B vssd1 vssd1 vccd1 vccd1 _5685_/C sky130_fd_sc_hd__nor2_2
X_8441_ input3/X _8441_/D vssd1 vssd1 vccd1 vccd1 _8441_/Q sky130_fd_sc_hd__dfxtp_1
X_4604_ _8455_/Q vssd1 vssd1 vccd1 vccd1 _5001_/A sky130_fd_sc_hd__inv_2
X_8372_ _8372_/A _8372_/B _8372_/C vssd1 vssd1 vccd1 vccd1 _8372_/Y sky130_fd_sc_hd__nand3_1
X_5584_ _5778_/A _5930_/A vssd1 vssd1 vccd1 vccd1 _6243_/B sky130_fd_sc_hd__or2_2
X_4535_ _4539_/C _4535_/B vssd1 vssd1 vccd1 vccd1 _8439_/D sky130_fd_sc_hd__nor2_1
X_7323_ _7323_/A _7323_/B vssd1 vssd1 vccd1 vccd1 _7324_/B sky130_fd_sc_hd__nor2_1
XFILLER_89_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7254_ _7352_/A _7254_/B vssd1 vssd1 vccd1 vccd1 _7349_/B sky130_fd_sc_hd__or2_1
X_4466_ _7518_/B _4466_/B _4715_/A _4713_/A vssd1 vssd1 vccd1 vccd1 _4591_/C sky130_fd_sc_hd__or4_1
XFILLER_89_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7185_ _7185_/A _7185_/B vssd1 vssd1 vccd1 vccd1 _7186_/B sky130_fd_sc_hd__nor2_1
X_4397_ _7554_/B vssd1 vssd1 vccd1 vccd1 _4638_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6205_ _6152_/A _6152_/B _5733_/B _6151_/S vssd1 vssd1 vccd1 vccd1 _6205_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_58_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6136_ _6030_/A _6030_/B _6135_/X vssd1 vssd1 vccd1 vccd1 _6143_/A sky130_fd_sc_hd__o21ai_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6067_ _6067_/A _6067_/B _6067_/C vssd1 vssd1 vccd1 vccd1 _6068_/B sky130_fd_sc_hd__nor3_1
XFILLER_45_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5018_ _5018_/A _5112_/A _5018_/C _5148_/C vssd1 vssd1 vccd1 vccd1 _5018_/X sky130_fd_sc_hd__or4_1
XFILLER_53_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6969_ _6969_/A _6969_/B _6969_/C vssd1 vssd1 vccd1 vccd1 _6970_/B sky130_fd_sc_hd__and3_1
XFILLER_41_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8708_ _8708_/A _4289_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[25] sky130_fd_sc_hd__ebufn_8
XFILLER_42_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4320_ _4320_/A vssd1 vssd1 vccd1 vccd1 _4320_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7941_ _7904_/A _7904_/B _7909_/A _7909_/B vssd1 vssd1 vccd1 vccd1 _8039_/A sky130_fd_sc_hd__a22oi_4
X_7872_ _8015_/A _7872_/B vssd1 vssd1 vccd1 vccd1 _8180_/B sky130_fd_sc_hd__xnor2_1
X_6823_ _6941_/A _6823_/B vssd1 vssd1 vccd1 vccd1 _6824_/B sky130_fd_sc_hd__xnor2_2
X_6754_ _7233_/B _7293_/A vssd1 vssd1 vccd1 vccd1 _6755_/B sky130_fd_sc_hd__or2_1
X_6685_ _7068_/B _6786_/B vssd1 vssd1 vccd1 vccd1 _6686_/C sky130_fd_sc_hd__nand2_1
X_5705_ _5705_/A _5984_/B vssd1 vssd1 vccd1 vccd1 _5706_/A sky130_fd_sc_hd__or2_1
XFILLER_31_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8424_ _8424_/A _8428_/B vssd1 vssd1 vccd1 vccd1 _8425_/B sky130_fd_sc_hd__nand2_1
X_5636_ _5720_/B _5635_/C _5635_/A vssd1 vssd1 vccd1 vccd1 _5636_/X sky130_fd_sc_hd__a21o_1
X_8355_ _8355_/A _8355_/B vssd1 vssd1 vccd1 vccd1 _8355_/Y sky130_fd_sc_hd__xnor2_1
X_5567_ _5578_/A _5567_/B vssd1 vssd1 vccd1 vccd1 _5586_/A sky130_fd_sc_hd__nand2_1
X_7306_ _7306_/A _6859_/A vssd1 vssd1 vccd1 vccd1 _7306_/X sky130_fd_sc_hd__or2b_1
X_8286_ _8286_/A _8296_/B vssd1 vssd1 vccd1 vccd1 _8297_/B sky130_fd_sc_hd__xnor2_1
XFILLER_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5498_ _5445_/A _5461_/A _5444_/B _5497_/Y vssd1 vssd1 vccd1 vccd1 _5499_/C sky130_fd_sc_hd__a31o_1
X_4518_ _8434_/Q _8433_/Q _8435_/Q vssd1 vssd1 vccd1 vccd1 _4527_/C sky130_fd_sc_hd__and3_1
X_4449_ _5121_/A vssd1 vssd1 vccd1 vccd1 _5016_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7237_ _7248_/A _7185_/A _7202_/Y _7070_/B vssd1 vssd1 vccd1 vccd1 _7244_/B sky130_fd_sc_hd__o22a_1
X_7168_ _7172_/A _7172_/B _7167_/X vssd1 vssd1 vccd1 vccd1 _7345_/C sky130_fd_sc_hd__a21boi_1
X_7099_ _7099_/A _7099_/B _7099_/C vssd1 vssd1 vccd1 vccd1 _7103_/A sky130_fd_sc_hd__nand3_1
X_6119_ _6216_/B _6119_/B vssd1 vssd1 vccd1 vccd1 _6122_/A sky130_fd_sc_hd__xnor2_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8674__90 vssd1 vssd1 vccd1 vccd1 _8674__90/HI _8783_/A sky130_fd_sc_hd__conb_1
XFILLER_76_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6470_ _7412_/A _6470_/B _6470_/C vssd1 vssd1 vccd1 vccd1 _6471_/A sky130_fd_sc_hd__and3_1
X_5421_ _5385_/A _5385_/B _5388_/B _5397_/X _5386_/X vssd1 vssd1 vccd1 vccd1 _5422_/B
+ sky130_fd_sc_hd__a311o_1
X_5352_ _5359_/B _5366_/A vssd1 vssd1 vccd1 vccd1 _5362_/A sky130_fd_sc_hd__or2b_1
X_8140_ _8140_/A _8140_/B vssd1 vssd1 vccd1 vccd1 _8141_/B sky130_fd_sc_hd__or2_1
X_4303_ _4327_/A vssd1 vssd1 vccd1 vccd1 _4308_/A sky130_fd_sc_hd__clkbuf_2
X_8071_ _8260_/A _8052_/B _8260_/B vssd1 vssd1 vccd1 vccd1 _8276_/B sky130_fd_sc_hd__a21o_1
X_7022_ _6954_/Y _7020_/X _7019_/Y _7019_/A vssd1 vssd1 vccd1 vccd1 _7022_/X sky130_fd_sc_hd__o211a_1
X_5283_ _8501_/Q _8502_/Q _5283_/C vssd1 vssd1 vccd1 vccd1 _5286_/B sky130_fd_sc_hd__and3_1
XINSDIODE2_9 _7351_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7924_ _8041_/A _7924_/B vssd1 vssd1 vccd1 vccd1 _7926_/C sky130_fd_sc_hd__xnor2_1
XFILLER_70_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7855_ _7855_/A _7855_/B vssd1 vssd1 vccd1 vccd1 _7856_/B sky130_fd_sc_hd__xnor2_1
XFILLER_36_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6806_ _6806_/A _6964_/B _6964_/C vssd1 vssd1 vccd1 vccd1 _6810_/B sky130_fd_sc_hd__or3_1
X_4998_ _5171_/A _4898_/A _4997_/X _4862_/B vssd1 vssd1 vccd1 vccd1 _4998_/X sky130_fd_sc_hd__o31a_1
XFILLER_51_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7786_ _7786_/A _7786_/B vssd1 vssd1 vccd1 vccd1 _7787_/B sky130_fd_sc_hd__and2_1
X_6737_ _6735_/Y _6736_/X _6643_/D vssd1 vssd1 vccd1 vccd1 _6802_/B sky130_fd_sc_hd__a21bo_1
X_6668_ _6569_/B _6580_/B _6569_/A vssd1 vssd1 vccd1 vccd1 _6669_/B sky130_fd_sc_hd__o21bai_2
X_6599_ _6736_/B vssd1 vssd1 vccd1 vccd1 _7038_/B sky130_fd_sc_hd__clkbuf_2
X_5619_ _5619_/A _5619_/B vssd1 vssd1 vccd1 vccd1 _5619_/X sky130_fd_sc_hd__xor2_1
X_8407_ _8401_/A _8401_/B _8399_/A vssd1 vssd1 vccd1 vccd1 _8414_/B sky130_fd_sc_hd__a21oi_1
X_8338_ _8284_/A _8339_/A vssd1 vssd1 vccd1 vccd1 _8338_/X sky130_fd_sc_hd__and2b_1
XFILLER_2_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8269_ _8269_/A _8269_/B vssd1 vssd1 vccd1 vccd1 _8281_/A sky130_fd_sc_hd__xnor2_1
XFILLER_93_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5970_ _5970_/A _5970_/B vssd1 vssd1 vccd1 vccd1 _5990_/A sky130_fd_sc_hd__nand2_1
X_4921_ _5090_/A _4921_/B vssd1 vssd1 vccd1 vccd1 _4921_/X sky130_fd_sc_hd__or2_2
X_4852_ _4944_/B _4796_/A _5011_/A vssd1 vssd1 vccd1 vccd1 _5036_/A sky130_fd_sc_hd__o21bai_4
X_7640_ _7546_/A _7768_/A _7526_/B _7639_/X vssd1 vssd1 vccd1 vccd1 _7657_/A sky130_fd_sc_hd__o31a_1
X_4783_ _5147_/A _4840_/A vssd1 vssd1 vccd1 vccd1 _5087_/A sky130_fd_sc_hd__or2_1
X_7571_ _7951_/A vssd1 vssd1 vccd1 vccd1 _7969_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_20_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6522_ _8566_/Q _8462_/Q vssd1 vssd1 vccd1 vccd1 _6522_/X sky130_fd_sc_hd__and2b_1
XFILLER_9_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6453_ _6452_/A _6459_/A _6452_/C vssd1 vssd1 vccd1 vccd1 _6453_/X sky130_fd_sc_hd__a21o_1
X_5404_ _5417_/A _5404_/B vssd1 vssd1 vccd1 vccd1 _5408_/B sky130_fd_sc_hd__xor2_2
X_6384_ _8545_/Q _6384_/B vssd1 vssd1 vccd1 vccd1 _6386_/A sky130_fd_sc_hd__and2_1
X_8123_ _8123_/A _8231_/B vssd1 vssd1 vccd1 vccd1 _8348_/A sky130_fd_sc_hd__xnor2_2
X_5335_ _5335_/A _8508_/Q vssd1 vssd1 vccd1 vccd1 _5336_/B sky130_fd_sc_hd__or2b_1
X_5266_ _5270_/C _5266_/B vssd1 vssd1 vccd1 vccd1 _8496_/D sky130_fd_sc_hd__nor2_1
X_8054_ _8054_/A _8054_/B vssd1 vssd1 vccd1 vccd1 _8248_/A sky130_fd_sc_hd__nor2_1
X_7005_ _7250_/A _7005_/B vssd1 vssd1 vccd1 vccd1 _7005_/X sky130_fd_sc_hd__or2_1
X_5197_ _8477_/Q _5205_/B vssd1 vssd1 vccd1 vccd1 _5197_/X sky130_fd_sc_hd__or2_1
XFILLER_28_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7907_ _8054_/B _7907_/B vssd1 vssd1 vccd1 vccd1 _7991_/A sky130_fd_sc_hd__nor2_2
XFILLER_70_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7838_ _7838_/A vssd1 vssd1 vccd1 vccd1 _7869_/A sky130_fd_sc_hd__inv_2
X_7769_ _7769_/A _7916_/A vssd1 vssd1 vccd1 vccd1 _8176_/A sky130_fd_sc_hd__nor2_2
XFILLER_59_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8644__60 vssd1 vssd1 vccd1 vccd1 _8644__60/HI _8753_/A sky130_fd_sc_hd__conb_1
XFILLER_93_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5120_ _5080_/A _5114_/X _5116_/X _5119_/X _4951_/A vssd1 vssd1 vccd1 vccd1 _5120_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5051_ _5051_/A _5116_/B vssd1 vssd1 vccd1 vccd1 _5058_/C sky130_fd_sc_hd__or2_1
XFILLER_38_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8741_ _8741_/A _4329_/Y vssd1 vssd1 vccd1 vccd1 io_out[26] sky130_fd_sc_hd__ebufn_8
XFILLER_65_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5953_ _5953_/A _5953_/B vssd1 vssd1 vccd1 vccd1 _6012_/B sky130_fd_sc_hd__xor2_1
X_4904_ _4960_/A _4955_/B _5041_/C _4996_/B vssd1 vssd1 vccd1 vccd1 _4904_/X sky130_fd_sc_hd__or4_1
X_5884_ _5884_/A _5914_/A vssd1 vssd1 vccd1 vccd1 _5885_/B sky130_fd_sc_hd__nor2_1
XFILLER_21_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4835_ _5104_/A vssd1 vssd1 vccd1 vccd1 _5019_/A sky130_fd_sc_hd__clkbuf_2
X_7623_ _7623_/A _7623_/B vssd1 vssd1 vccd1 vccd1 _7624_/B sky130_fd_sc_hd__xor2_1
X_4766_ _8465_/Q _4766_/B _4766_/C vssd1 vssd1 vccd1 vccd1 _4817_/A sky130_fd_sc_hd__or3_4
XFILLER_21_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7554_ _8583_/Q _7554_/B vssd1 vssd1 vccd1 vccd1 _7556_/A sky130_fd_sc_hd__and2b_1
X_6505_ _6505_/A _6505_/B vssd1 vssd1 vccd1 vccd1 _6509_/A sky130_fd_sc_hd__xor2_2
X_4697_ _4698_/B _4698_/C _4698_/A vssd1 vssd1 vccd1 vccd1 _4699_/B sky130_fd_sc_hd__a21o_1
X_7485_ _8426_/A _7485_/B vssd1 vssd1 vccd1 vccd1 _7485_/Y sky130_fd_sc_hd__nor2_1
X_6436_ _6434_/Y _6436_/B vssd1 vssd1 vccd1 vccd1 _6436_/X sky130_fd_sc_hd__and2b_1
X_6367_ _8539_/Q _6366_/B _6348_/X vssd1 vssd1 vccd1 vccd1 _6368_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8106_ _7984_/A _7925_/B _8123_/A _8096_/X vssd1 vssd1 vccd1 vccd1 _8107_/B sky130_fd_sc_hd__a31oi_1
X_5318_ _5360_/A _5366_/A _5317_/X _8515_/Q vssd1 vssd1 vccd1 vccd1 _5318_/Y sky130_fd_sc_hd__a31oi_1
X_6298_ _6294_/A _6297_/X _6298_/S vssd1 vssd1 vccd1 vccd1 _6298_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5249_ _5249_/A vssd1 vssd1 vccd1 vccd1 _8491_/D sky130_fd_sc_hd__clkbuf_1
X_8037_ _8037_/A _8037_/B vssd1 vssd1 vccd1 vccd1 _8038_/B sky130_fd_sc_hd__nand2_1
XFILLER_56_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4620_ _4620_/A vssd1 vssd1 vccd1 vccd1 _4640_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4551_ _4551_/A vssd1 vssd1 vccd1 vccd1 _8444_/D sky130_fd_sc_hd__clkbuf_1
X_7270_ _7270_/A _7270_/B vssd1 vssd1 vccd1 vccd1 _7356_/A sky130_fd_sc_hd__nand2_2
X_4482_ _4495_/B vssd1 vssd1 vccd1 vccd1 _4491_/B sky130_fd_sc_hd__clkbuf_1
X_6221_ _6221_/A _6221_/B vssd1 vssd1 vccd1 vccd1 _6222_/B sky130_fd_sc_hd__xnor2_1
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6152_ _6152_/A _6152_/B vssd1 vssd1 vccd1 vccd1 _6156_/A sky130_fd_sc_hd__xor2_1
X_5103_ _5171_/A _5132_/C _5100_/X _5102_/X vssd1 vssd1 vccd1 vccd1 _5103_/X sky130_fd_sc_hd__o31a_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6083_ _6090_/D _6083_/B vssd1 vssd1 vccd1 vccd1 _6086_/A sky130_fd_sc_hd__nand2_1
X_5034_ _5109_/C _5027_/X _5028_/X _5033_/X vssd1 vssd1 vccd1 vccd1 _5034_/X sky130_fd_sc_hd__o31a_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6985_ _6985_/A _6985_/B vssd1 vssd1 vccd1 vccd1 _7062_/A sky130_fd_sc_hd__xor2_2
XFILLER_41_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8724_ _8724_/A _4308_/Y vssd1 vssd1 vccd1 vccd1 io_out[9] sky130_fd_sc_hd__ebufn_8
XFILLER_15_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5936_ _6008_/A _5936_/B vssd1 vssd1 vccd1 vccd1 _5955_/A sky130_fd_sc_hd__nand2_1
XFILLER_80_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5867_ _5924_/A _5867_/B vssd1 vssd1 vccd1 vccd1 _5868_/B sky130_fd_sc_hd__and2_1
XFILLER_21_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7606_ _7606_/A _7606_/B vssd1 vssd1 vccd1 vccd1 _7607_/B sky130_fd_sc_hd__xor2_1
X_4818_ _4944_/A _4818_/B vssd1 vssd1 vccd1 vccd1 _5080_/B sky130_fd_sc_hd__nor2_2
X_5798_ _5861_/C vssd1 vssd1 vccd1 vccd1 _6126_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_31_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8586_ input3/X _8586_/D vssd1 vssd1 vccd1 vccd1 _8586_/Q sky130_fd_sc_hd__dfxtp_1
X_4749_ _4749_/A vssd1 vssd1 vccd1 vccd1 _4750_/A sky130_fd_sc_hd__inv_2
X_7537_ _7537_/A _7537_/B vssd1 vssd1 vccd1 vccd1 _8367_/A sky130_fd_sc_hd__nand2_2
X_7468_ _7466_/X _7467_/X _7399_/B vssd1 vssd1 vccd1 vccd1 _7468_/Y sky130_fd_sc_hd__o21ai_1
X_6419_ _6433_/A _8550_/Q _6450_/B _6439_/A _6445_/A vssd1 vssd1 vccd1 vccd1 _6419_/X
+ sky130_fd_sc_hd__a2111o_1
X_7399_ _8565_/Q _7399_/B _7410_/B vssd1 vssd1 vccd1 vccd1 _7399_/X sky130_fd_sc_hd__and3_1
XFILLER_88_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8614__30 vssd1 vssd1 vccd1 vccd1 _8614__30/HI _8709_/A sky130_fd_sc_hd__conb_1
XFILLER_29_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6770_ _6771_/A _6771_/B vssd1 vssd1 vccd1 vccd1 _6828_/A sky130_fd_sc_hd__nor2_2
XFILLER_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5721_ _5620_/A _5721_/B vssd1 vssd1 vccd1 vccd1 _5736_/A sky130_fd_sc_hd__and2b_1
XFILLER_50_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5652_ _5408_/B _5800_/B _5900_/B vssd1 vssd1 vccd1 vccd1 _5653_/B sky130_fd_sc_hd__a21oi_1
X_8440_ input3/X _8440_/D vssd1 vssd1 vccd1 vccd1 _8440_/Q sky130_fd_sc_hd__dfxtp_1
X_4603_ _4592_/A _4663_/A _4619_/B _4602_/X vssd1 vssd1 vccd1 vccd1 _8454_/D sky130_fd_sc_hd__o211a_1
X_8371_ _8371_/A _8376_/B vssd1 vssd1 vccd1 vccd1 _8372_/C sky130_fd_sc_hd__nand2_1
X_5583_ _5932_/A _5583_/B vssd1 vssd1 vccd1 vccd1 _5930_/A sky130_fd_sc_hd__nand2_1
X_7322_ _6783_/A _6783_/B _7321_/X vssd1 vssd1 vccd1 vccd1 _7324_/A sky130_fd_sc_hd__o21a_1
XFILLER_7_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4534_ _8439_/Q _4532_/A _4524_/X vssd1 vssd1 vccd1 vccd1 _4535_/B sky130_fd_sc_hd__o21ai_1
X_7253_ _7253_/A _7253_/B _7359_/A vssd1 vssd1 vccd1 vccd1 _7254_/B sky130_fd_sc_hd__nor3_1
X_4465_ _8473_/Q vssd1 vssd1 vccd1 vccd1 _5526_/B sky130_fd_sc_hd__clkbuf_2
X_7184_ _7248_/B _7184_/B _7184_/C vssd1 vssd1 vccd1 vccd1 _7185_/A sky130_fd_sc_hd__and3_2
X_4396_ _8459_/Q vssd1 vssd1 vccd1 vccd1 _7554_/B sky130_fd_sc_hd__clkbuf_4
X_6204_ _6204_/A _6204_/B vssd1 vssd1 vccd1 vccd1 _6207_/A sky130_fd_sc_hd__xnor2_1
X_6135_ _6135_/A _6135_/B vssd1 vssd1 vccd1 vccd1 _6135_/X sky130_fd_sc_hd__or2_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6066_ _6078_/A _6078_/B _6078_/C vssd1 vssd1 vccd1 vccd1 _6079_/A sky130_fd_sc_hd__o21a_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5017_ _5132_/C _5009_/X _5015_/X _5016_/X vssd1 vssd1 vccd1 vccd1 _5017_/X sky130_fd_sc_hd__o22a_1
XFILLER_85_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8707_ _8707_/A _4288_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[24] sky130_fd_sc_hd__ebufn_8
X_6968_ _6972_/A vssd1 vssd1 vccd1 vccd1 _6969_/A sky130_fd_sc_hd__inv_2
XFILLER_53_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6899_ _6899_/A _6899_/B _6899_/C vssd1 vssd1 vccd1 vccd1 _6924_/A sky130_fd_sc_hd__nand3_4
X_5919_ _6184_/A _5902_/X _5857_/Y vssd1 vssd1 vccd1 vccd1 _5921_/B sky130_fd_sc_hd__a21o_1
XFILLER_42_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8569_ input3/X _8569_/D vssd1 vssd1 vccd1 vccd1 _8569_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7940_ _7935_/A _7935_/B _7939_/Y vssd1 vssd1 vccd1 vccd1 _7996_/A sky130_fd_sc_hd__o21a_1
XFILLER_82_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7871_ _7933_/B _7871_/B vssd1 vssd1 vccd1 vccd1 _8015_/A sky130_fd_sc_hd__nand2_1
X_6822_ _6822_/A _6822_/B vssd1 vssd1 vccd1 vccd1 _6824_/A sky130_fd_sc_hd__xnor2_2
XFILLER_23_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6753_ _6842_/B vssd1 vssd1 vccd1 vccd1 _7293_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_50_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6684_ _7001_/B _7184_/B vssd1 vssd1 vccd1 vccd1 _7005_/B sky130_fd_sc_hd__nand2_2
X_5704_ _5855_/B vssd1 vssd1 vccd1 vccd1 _5984_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_31_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5635_ _5635_/A _5720_/B _5635_/C vssd1 vssd1 vccd1 vccd1 _5718_/A sky130_fd_sc_hd__nand3_1
X_8423_ _8423_/A _8423_/B vssd1 vssd1 vccd1 vccd1 _8428_/B sky130_fd_sc_hd__or2_1
X_5566_ _6244_/A _5410_/A _5980_/C _5565_/Y _5413_/X vssd1 vssd1 vccd1 vccd1 _5567_/B
+ sky130_fd_sc_hd__a32o_1
X_8354_ _8355_/A _8355_/B _8204_/A vssd1 vssd1 vccd1 vccd1 _8354_/Y sky130_fd_sc_hd__a21oi_1
X_7305_ _6660_/A _6647_/B _6824_/A _7304_/Y vssd1 vssd1 vccd1 vccd1 _7308_/A sky130_fd_sc_hd__a31o_1
X_8285_ _8285_/A _8285_/B vssd1 vssd1 vccd1 vccd1 _8296_/B sky130_fd_sc_hd__xnor2_1
X_5497_ _5497_/A _5497_/B vssd1 vssd1 vccd1 vccd1 _5497_/Y sky130_fd_sc_hd__nand2_1
X_4517_ _4517_/A vssd1 vssd1 vccd1 vccd1 _8434_/D sky130_fd_sc_hd__clkbuf_1
X_4448_ _8456_/Q vssd1 vssd1 vccd1 vccd1 _5121_/A sky130_fd_sc_hd__clkbuf_2
X_7236_ _7247_/A _7236_/B vssd1 vssd1 vccd1 vccd1 _7244_/A sky130_fd_sc_hd__xnor2_1
X_7167_ _7167_/A _7166_/B vssd1 vssd1 vccd1 vccd1 _7167_/X sky130_fd_sc_hd__or2b_1
XFILLER_86_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4379_ _4381_/A vssd1 vssd1 vccd1 vccd1 _4379_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7098_ _7098_/A _7098_/B _7264_/A vssd1 vssd1 vccd1 vccd1 _7268_/B sky130_fd_sc_hd__or3_1
XFILLER_85_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6118_ _6118_/A _6118_/B vssd1 vssd1 vccd1 vccd1 _6119_/B sky130_fd_sc_hd__xnor2_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6049_ _5964_/Y _6050_/A vssd1 vssd1 vccd1 vccd1 _6169_/A sky130_fd_sc_hd__nand2b_1
XFILLER_37_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5420_ _5420_/A _5419_/Y vssd1 vssd1 vccd1 vccd1 _5532_/A sky130_fd_sc_hd__nor2b_4
X_5351_ _5345_/B _5326_/B _5349_/Y _5350_/X _4668_/X vssd1 vssd1 vccd1 vccd1 _8512_/D
+ sky130_fd_sc_hd__o221a_1
X_4302_ input1/X vssd1 vssd1 vccd1 vccd1 _4327_/A sky130_fd_sc_hd__clkbuf_2
X_5282_ _5282_/A _5282_/B vssd1 vssd1 vccd1 vccd1 _8501_/D sky130_fd_sc_hd__nor2_1
X_8070_ _8070_/A _8155_/B vssd1 vssd1 vccd1 vccd1 _8072_/A sky130_fd_sc_hd__xnor2_1
X_7021_ _7019_/A _7019_/Y _7020_/X _6954_/Y vssd1 vssd1 vccd1 vccd1 _7021_/Y sky130_fd_sc_hd__a211oi_4
XFILLER_68_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7923_ _7808_/A _8249_/A _7922_/Y vssd1 vssd1 vccd1 vccd1 _7924_/B sky130_fd_sc_hd__o21a_1
XFILLER_82_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7854_ _8069_/A _7854_/B vssd1 vssd1 vccd1 vccd1 _7855_/B sky130_fd_sc_hd__nor2_1
XFILLER_36_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6805_ _6643_/D _6739_/B _6736_/X vssd1 vssd1 vccd1 vccd1 _6836_/A sky130_fd_sc_hd__o21ai_1
X_7785_ _7786_/A _7786_/B vssd1 vssd1 vccd1 vccd1 _8198_/A sky130_fd_sc_hd__nor2_1
X_4997_ _4584_/A _4992_/X _4996_/X vssd1 vssd1 vccd1 vccd1 _4997_/X sky130_fd_sc_hd__o21a_1
X_6736_ _6736_/A _6736_/B vssd1 vssd1 vccd1 vccd1 _6736_/X sky130_fd_sc_hd__or2_1
XFILLER_23_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6667_ _7118_/A _6721_/A vssd1 vssd1 vccd1 vccd1 _7079_/A sky130_fd_sc_hd__xnor2_4
X_6598_ _6964_/C vssd1 vssd1 vccd1 vccd1 _6736_/B sky130_fd_sc_hd__clkbuf_2
X_5618_ _5618_/A _5627_/A vssd1 vssd1 vccd1 vccd1 _5619_/B sky130_fd_sc_hd__xnor2_1
X_8406_ _8415_/A _8406_/B vssd1 vssd1 vccd1 vccd1 _8408_/A sky130_fd_sc_hd__or2_1
X_8337_ _8337_/A _8337_/B vssd1 vssd1 vccd1 vccd1 _8342_/A sky130_fd_sc_hd__xnor2_1
XFILLER_3_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5549_ _5537_/B _5427_/Y _5539_/B vssd1 vssd1 vccd1 vccd1 _5551_/B sky130_fd_sc_hd__o21ai_1
X_8268_ _8054_/B _8142_/B _8141_/A vssd1 vssd1 vccd1 vccd1 _8269_/B sky130_fd_sc_hd__o21a_1
X_7219_ _7219_/A _7219_/B vssd1 vssd1 vccd1 vccd1 _7234_/A sky130_fd_sc_hd__xnor2_2
XFILLER_59_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8199_ _8199_/A _8199_/B vssd1 vssd1 vccd1 vccd1 _8211_/B sky130_fd_sc_hd__xnor2_1
XFILLER_86_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4920_ _4955_/A _5064_/C vssd1 vssd1 vccd1 vccd1 _4920_/X sky130_fd_sc_hd__or2_1
XFILLER_64_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4851_ _5136_/B vssd1 vssd1 vccd1 vccd1 _5132_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_33_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4782_ _4899_/A _4782_/B vssd1 vssd1 vccd1 vccd1 _4840_/A sky130_fd_sc_hd__nor2_1
XFILLER_60_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7570_ _7888_/A vssd1 vssd1 vccd1 vccd1 _7951_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6521_ _6521_/A _6521_/B vssd1 vssd1 vccd1 vccd1 _6521_/X sky130_fd_sc_hd__and2_1
XFILLER_20_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6452_ _6452_/A _6459_/A _6452_/C vssd1 vssd1 vccd1 vccd1 _6466_/A sky130_fd_sc_hd__nand3_1
X_5403_ _5800_/A vssd1 vssd1 vccd1 vccd1 _5694_/A sky130_fd_sc_hd__clkbuf_2
X_6383_ _6383_/A vssd1 vssd1 vccd1 vccd1 _8544_/D sky130_fd_sc_hd__clkbuf_1
X_8122_ _7813_/A _7984_/C _8249_/B vssd1 vssd1 vccd1 vccd1 _8231_/B sky130_fd_sc_hd__mux2_1
X_5334_ _8508_/Q _5335_/A vssd1 vssd1 vccd1 vccd1 _5336_/A sky130_fd_sc_hd__or2b_1
X_5265_ _8496_/Q _5263_/B _5264_/X vssd1 vssd1 vccd1 vccd1 _5266_/B sky130_fd_sc_hd__o21ai_1
X_8053_ _8366_/B _8053_/B _8053_/C vssd1 vssd1 vccd1 vccd1 _8323_/A sky130_fd_sc_hd__and3_1
X_5196_ _8518_/Q _5188_/X _5195_/X _6426_/A vssd1 vssd1 vccd1 vccd1 _8476_/D sky130_fd_sc_hd__o211a_1
X_7004_ _7250_/A _7005_/B _7003_/X vssd1 vssd1 vccd1 vccd1 _7148_/B sky130_fd_sc_hd__o21ai_4
XFILLER_18_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7906_ _7747_/A _8054_/B _7866_/B _7865_/A vssd1 vssd1 vccd1 vccd1 _7907_/B sky130_fd_sc_hd__o31a_1
XFILLER_51_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7837_ _7837_/A _7837_/B vssd1 vssd1 vccd1 vccd1 _7873_/B sky130_fd_sc_hd__nand2_2
XFILLER_36_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7768_ _7768_/A _7978_/B vssd1 vssd1 vccd1 vccd1 _7916_/A sky130_fd_sc_hd__or2_1
X_6719_ _6938_/A _6938_/B _6718_/X vssd1 vssd1 vccd1 vccd1 _6937_/B sky130_fd_sc_hd__o21ai_1
XFILLER_50_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7699_ _8054_/A _7699_/B vssd1 vssd1 vccd1 vccd1 _8052_/B sky130_fd_sc_hd__nand2_1
XFILLER_50_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5050_ _5050_/A _5160_/A _5050_/C vssd1 vssd1 vccd1 vccd1 _5050_/X sky130_fd_sc_hd__or3_1
XFILLER_69_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8740_ _8740_/A _4328_/Y vssd1 vssd1 vccd1 vccd1 io_out[25] sky130_fd_sc_hd__ebufn_8
XFILLER_65_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5952_ _5952_/A _6037_/B vssd1 vssd1 vccd1 vccd1 _5953_/B sky130_fd_sc_hd__xnor2_1
X_4903_ _5071_/A _5055_/B _5071_/C vssd1 vssd1 vccd1 vccd1 _4996_/B sky130_fd_sc_hd__or3_2
XFILLER_80_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5883_ _6244_/B _5689_/A _5992_/A vssd1 vssd1 vccd1 vccd1 _5884_/A sky130_fd_sc_hd__a21oi_1
XFILLER_21_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4834_ _4713_/A _4609_/A _4592_/A _4827_/X _4833_/X vssd1 vssd1 vccd1 vccd1 _4834_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_21_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7622_ _7744_/A _7744_/B vssd1 vssd1 vccd1 vccd1 _7623_/B sky130_fd_sc_hd__xor2_1
X_4765_ _4765_/A _4765_/B vssd1 vssd1 vccd1 vccd1 _4943_/B sky130_fd_sc_hd__nor2_2
X_7553_ _7553_/A _7553_/B vssd1 vssd1 vccd1 vccd1 _7576_/A sky130_fd_sc_hd__or2_1
X_6504_ _7202_/A _6508_/C _6585_/C vssd1 vssd1 vccd1 vccd1 _6505_/B sky130_fd_sc_hd__o21a_1
X_4696_ _4696_/A vssd1 vssd1 vccd1 vccd1 _8470_/D sky130_fd_sc_hd__clkbuf_1
X_7484_ _7484_/A _7484_/B vssd1 vssd1 vccd1 vccd1 _7485_/B sky130_fd_sc_hd__xnor2_1
X_6435_ _6435_/A _6435_/B vssd1 vssd1 vccd1 vccd1 _6436_/B sky130_fd_sc_hd__nand2_1
XFILLER_20_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6366_ _8539_/Q _6366_/B vssd1 vssd1 vccd1 vccd1 _6371_/C sky130_fd_sc_hd__and2_1
XFILLER_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8105_ _8105_/A _8105_/B vssd1 vssd1 vccd1 vccd1 _8123_/A sky130_fd_sc_hd__nor2_2
X_5317_ _5335_/A _8509_/Q _5345_/B _5339_/B vssd1 vssd1 vccd1 vccd1 _5317_/X sky130_fd_sc_hd__a211o_1
X_8036_ _8086_/A _8086_/B vssd1 vssd1 vccd1 vccd1 _8038_/A sky130_fd_sc_hd__xor2_1
XFILLER_29_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6297_ _6286_/B _6297_/B vssd1 vssd1 vccd1 vccd1 _6297_/X sky130_fd_sc_hd__and2b_1
X_5248_ _5253_/C _5248_/B _5291_/A vssd1 vssd1 vccd1 vccd1 _5249_/A sky130_fd_sc_hd__and3b_1
X_5179_ _5179_/A _5179_/B vssd1 vssd1 vccd1 vccd1 _5179_/Y sky130_fd_sc_hd__nand2_1
XFILLER_29_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4550_ _4552_/B _4568_/B _4550_/C vssd1 vssd1 vccd1 vccd1 _4551_/A sky130_fd_sc_hd__and3b_1
X_4481_ _4481_/A vssd1 vssd1 vccd1 vccd1 _8736_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6220_ _6220_/A _6220_/B vssd1 vssd1 vccd1 vccd1 _6221_/B sky130_fd_sc_hd__xnor2_1
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6151_ _5778_/X _6150_/Y _6151_/S vssd1 vssd1 vccd1 vccd1 _6152_/B sky130_fd_sc_hd__mux2_1
X_5102_ _5102_/A _5107_/C _5104_/B _5102_/D vssd1 vssd1 vccd1 vccd1 _5102_/X sky130_fd_sc_hd__or4_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6082_ _6082_/A _6082_/B _6083_/B vssd1 vssd1 vccd1 vccd1 _6238_/A sky130_fd_sc_hd__and3_1
X_5033_ _5102_/A _5099_/B _5033_/C _5033_/D vssd1 vssd1 vccd1 vccd1 _5033_/X sky130_fd_sc_hd__or4_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6984_ _6985_/A _6985_/B vssd1 vssd1 vccd1 vccd1 _6984_/X sky130_fd_sc_hd__or2_2
XFILLER_53_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8723_ _8723_/A _4307_/Y vssd1 vssd1 vccd1 vccd1 io_out[8] sky130_fd_sc_hd__ebufn_8
XFILLER_15_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5935_ _5935_/A _5935_/B vssd1 vssd1 vccd1 vccd1 _5936_/B sky130_fd_sc_hd__or2_1
X_5866_ _5866_/A _6129_/A vssd1 vssd1 vccd1 vccd1 _5867_/B sky130_fd_sc_hd__or2_1
X_4817_ _4817_/A _4953_/B vssd1 vssd1 vccd1 vccd1 _4938_/A sky130_fd_sc_hd__nor2_2
XFILLER_21_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7605_ _7888_/A _7725_/C vssd1 vssd1 vccd1 vccd1 _7744_/A sky130_fd_sc_hd__nor2_2
X_5797_ _5978_/B vssd1 vssd1 vccd1 vccd1 _5861_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_21_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8585_ input3/X _8585_/D vssd1 vssd1 vccd1 vccd1 _8585_/Q sky130_fd_sc_hd__dfxtp_1
X_4748_ _4735_/A _4748_/B _4759_/B _4748_/D vssd1 vssd1 vccd1 vccd1 _4749_/A sky130_fd_sc_hd__and4b_1
X_7536_ _8023_/A _7528_/C _7804_/A vssd1 vssd1 vccd1 vccd1 _7549_/B sky130_fd_sc_hd__o21a_1
X_4679_ _4671_/B _4808_/A _4677_/X _5207_/A _4780_/A vssd1 vssd1 vccd1 vccd1 _4680_/B
+ sky130_fd_sc_hd__a32o_1
X_7467_ _7459_/A _7461_/B _7459_/B vssd1 vssd1 vccd1 vccd1 _7467_/X sky130_fd_sc_hd__o21ba_1
X_6418_ _8553_/Q vssd1 vssd1 vccd1 vccd1 _6445_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7398_ _7398_/A _7398_/B vssd1 vssd1 vccd1 vccd1 _7398_/Y sky130_fd_sc_hd__nand2_1
X_6349_ _6351_/A _6351_/C _6348_/X vssd1 vssd1 vccd1 vccd1 _6350_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8019_ _7996_/A _8019_/B vssd1 vssd1 vccd1 vccd1 _8019_/X sky130_fd_sc_hd__and2b_1
XFILLER_56_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5720_ _5633_/A _5720_/B vssd1 vssd1 vccd1 vccd1 _5744_/A sky130_fd_sc_hd__and2b_1
XFILLER_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5651_ _5651_/A _5855_/B vssd1 vssd1 vccd1 vccd1 _5900_/B sky130_fd_sc_hd__nor2_2
XFILLER_30_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4602_ _4657_/B vssd1 vssd1 vccd1 vccd1 _4602_/X sky130_fd_sc_hd__clkbuf_2
X_8370_ _8370_/A _8370_/B vssd1 vssd1 vccd1 vccd1 _8376_/B sky130_fd_sc_hd__xnor2_1
X_5582_ _5828_/A _5738_/A vssd1 vssd1 vccd1 vccd1 _5583_/B sky130_fd_sc_hd__nand2_1
X_7321_ _7321_/A _7321_/B vssd1 vssd1 vccd1 vccd1 _7321_/X sky130_fd_sc_hd__or2_1
X_4533_ _8438_/Q _8439_/Q _4533_/C vssd1 vssd1 vccd1 vccd1 _4539_/C sky130_fd_sc_hd__and3_1
X_7252_ _7358_/A _7358_/B vssd1 vssd1 vccd1 vccd1 _7359_/A sky130_fd_sc_hd__or2_1
XFILLER_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4464_ _4713_/A _4464_/B _4464_/C _4805_/A vssd1 vssd1 vccd1 vccd1 _4470_/C sky130_fd_sc_hd__or4_1
X_6203_ _5948_/A _6151_/S _6150_/Y vssd1 vssd1 vccd1 vccd1 _6204_/B sky130_fd_sc_hd__o21a_1
X_4395_ _8460_/Q vssd1 vssd1 vccd1 vccd1 _7575_/B sky130_fd_sc_hd__clkbuf_4
X_7183_ _7183_/A _7202_/B vssd1 vssd1 vccd1 vccd1 _7184_/C sky130_fd_sc_hd__nor2_1
X_6134_ _6134_/A _6134_/B vssd1 vssd1 vccd1 vccd1 _6163_/A sky130_fd_sc_hd__xnor2_1
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6065_ _6065_/A _6065_/B vssd1 vssd1 vccd1 vccd1 _6078_/C sky130_fd_sc_hd__xor2_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5016_ _5016_/A _5031_/B _5095_/C vssd1 vssd1 vccd1 vccd1 _5016_/X sky130_fd_sc_hd__or3_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6967_ _6977_/A _7044_/A _7044_/B _7034_/S vssd1 vssd1 vccd1 vccd1 _6967_/X sky130_fd_sc_hd__a31o_1
XFILLER_14_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8706_ _8706_/A _4287_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[23] sky130_fd_sc_hd__ebufn_8
XFILLER_53_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5918_ _5918_/A _5992_/A _5918_/C vssd1 vssd1 vccd1 vccd1 _6006_/A sky130_fd_sc_hd__and3_1
XFILLER_41_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6898_ _6896_/A _6896_/B _6896_/C vssd1 vssd1 vccd1 vccd1 _6899_/C sky130_fd_sc_hd__a21o_1
X_5849_ _5776_/A _5776_/B _5780_/B _5781_/B _5781_/A vssd1 vssd1 vccd1 vccd1 _5851_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_42_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8568_ input3/X _8568_/D vssd1 vssd1 vccd1 vccd1 _8568_/Q sky130_fd_sc_hd__dfxtp_1
X_7519_ _7517_/X _7542_/A vssd1 vssd1 vccd1 vccd1 _7520_/B sky130_fd_sc_hd__and2b_1
X_8499_ input3/X _8499_/D vssd1 vssd1 vccd1 vccd1 _8499_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7870_ _7873_/B _7870_/B vssd1 vssd1 vccd1 vccd1 _8180_/A sky130_fd_sc_hd__xnor2_1
X_6821_ _7286_/A _7286_/B vssd1 vssd1 vccd1 vccd1 _6822_/B sky130_fd_sc_hd__xor2_2
XFILLER_23_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6752_ _7032_/A vssd1 vssd1 vccd1 vccd1 _7233_/B sky130_fd_sc_hd__buf_2
XFILLER_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6683_ _6683_/A _6683_/B vssd1 vssd1 vccd1 vccd1 _7184_/B sky130_fd_sc_hd__nor2_1
X_5703_ _5703_/A _5800_/B vssd1 vssd1 vccd1 vccd1 _6183_/S sky130_fd_sc_hd__nand2_2
X_5634_ _5633_/A _5633_/B _5632_/X vssd1 vssd1 vccd1 vccd1 _5635_/C sky130_fd_sc_hd__o21bai_1
X_8422_ _8423_/A _8423_/B vssd1 vssd1 vccd1 vccd1 _8424_/A sky130_fd_sc_hd__nand2_1
X_8353_ _8353_/A _8353_/B vssd1 vssd1 vccd1 vccd1 _8385_/B sky130_fd_sc_hd__xnor2_4
X_7304_ _6660_/A _6702_/A _6824_/A _6824_/B vssd1 vssd1 vccd1 vccd1 _7304_/Y sky130_fd_sc_hd__a211oi_1
X_5565_ _5565_/A _5565_/B vssd1 vssd1 vccd1 vccd1 _5565_/Y sky130_fd_sc_hd__nand2_1
X_8284_ _8284_/A _8339_/A vssd1 vssd1 vccd1 vccd1 _8285_/B sky130_fd_sc_hd__xnor2_1
XFILLER_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5496_ _5494_/X _5496_/B vssd1 vssd1 vccd1 vccd1 _5499_/B sky130_fd_sc_hd__and2b_1
X_4516_ _4516_/A _4575_/A _4516_/C vssd1 vssd1 vccd1 vccd1 _4517_/A sky130_fd_sc_hd__and3_1
X_4447_ _6482_/B vssd1 vssd1 vccd1 vccd1 _4624_/A sky130_fd_sc_hd__clkbuf_2
X_7235_ _7247_/A _7236_/B vssd1 vssd1 vccd1 vccd1 _7239_/A sky130_fd_sc_hd__and2b_1
X_7166_ _7167_/A _7166_/B vssd1 vssd1 vccd1 vccd1 _7172_/B sky130_fd_sc_hd__xnor2_1
X_4378_ _4381_/A vssd1 vssd1 vccd1 vccd1 _4378_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6117_ _6117_/A _6117_/B vssd1 vssd1 vccd1 vccd1 _6118_/B sky130_fd_sc_hd__xor2_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7097_ _7030_/X _7097_/B vssd1 vssd1 vccd1 vccd1 _7268_/A sky130_fd_sc_hd__and2b_1
XFILLER_85_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6048_ _6048_/A _6048_/B vssd1 vssd1 vccd1 vccd1 _6050_/A sky130_fd_sc_hd__xor2_1
XFILLER_85_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7999_ _7808_/A _8249_/A _7998_/X vssd1 vssd1 vccd1 vccd1 _8022_/B sky130_fd_sc_hd__o21ai_1
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5350_ _5349_/A _5349_/B _5368_/B vssd1 vssd1 vccd1 vccd1 _5350_/X sky130_fd_sc_hd__a21o_1
X_4301_ _4301_/A vssd1 vssd1 vccd1 vccd1 _4301_/Y sky130_fd_sc_hd__inv_2
X_5281_ _8501_/Q _5283_/C _5264_/X vssd1 vssd1 vccd1 vccd1 _5282_/B sky130_fd_sc_hd__o21ai_1
XFILLER_87_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7020_ _6954_/A _6954_/B _6954_/C vssd1 vssd1 vccd1 vccd1 _7020_/X sky130_fd_sc_hd__o21a_1
X_8665__81 vssd1 vssd1 vccd1 vccd1 _8665__81/HI _8774_/A sky130_fd_sc_hd__conb_1
XFILLER_67_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7922_ _8041_/C _8025_/A vssd1 vssd1 vccd1 vccd1 _7922_/Y sky130_fd_sc_hd__nand2_1
XFILLER_82_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7853_ _7962_/A _7945_/A vssd1 vssd1 vccd1 vccd1 _7854_/B sky130_fd_sc_hd__and2_1
XFILLER_23_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4996_ _4996_/A _4996_/B _4996_/C vssd1 vssd1 vccd1 vccd1 _4996_/X sky130_fd_sc_hd__or3_1
X_6804_ _6804_/A _6804_/B vssd1 vssd1 vccd1 vccd1 _6839_/A sky130_fd_sc_hd__nand2_1
XFILLER_51_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7784_ _7782_/Y _7783_/X _7656_/B _7665_/A vssd1 vssd1 vccd1 vccd1 _7786_/B sky130_fd_sc_hd__o31a_1
X_6735_ _7175_/B _7032_/C _6842_/B vssd1 vssd1 vccd1 vccd1 _6735_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_51_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6666_ _6926_/A vssd1 vssd1 vccd1 vccd1 _7118_/A sky130_fd_sc_hd__buf_4
X_6597_ _6597_/A _6597_/B vssd1 vssd1 vccd1 vccd1 _6964_/C sky130_fd_sc_hd__xnor2_2
X_5617_ _5774_/A _5767_/B vssd1 vssd1 vccd1 vccd1 _5627_/A sky130_fd_sc_hd__or2_1
X_8405_ _8405_/A _8423_/B vssd1 vssd1 vccd1 vccd1 _8406_/B sky130_fd_sc_hd__nor2_1
X_8336_ _8336_/A _8336_/B vssd1 vssd1 vccd1 vccd1 _8337_/B sky130_fd_sc_hd__xnor2_1
X_5548_ _5548_/A _5548_/B vssd1 vssd1 vccd1 vccd1 _5551_/A sky130_fd_sc_hd__nand2_1
X_8267_ _8267_/A _8267_/B vssd1 vssd1 vccd1 vccd1 _8269_/A sky130_fd_sc_hd__nand2_1
X_7218_ _7218_/A _7218_/B vssd1 vssd1 vccd1 vccd1 _7256_/A sky130_fd_sc_hd__xor2_1
X_5479_ _5938_/A _5828_/A vssd1 vssd1 vccd1 vccd1 _5602_/A sky130_fd_sc_hd__or2_1
X_8198_ _8198_/A _8198_/B vssd1 vssd1 vccd1 vccd1 _8199_/A sky130_fd_sc_hd__nand2_1
X_7149_ _7149_/A _7149_/B vssd1 vssd1 vccd1 vccd1 _7181_/B sky130_fd_sc_hd__xnor2_1
XFILLER_48_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4850_ _5064_/B vssd1 vssd1 vccd1 vccd1 _5136_/B sky130_fd_sc_hd__clkbuf_2
X_4781_ _4899_/A _4875_/B _4994_/B vssd1 vssd1 vccd1 vccd1 _5147_/A sky130_fd_sc_hd__o21ai_4
X_6520_ _6999_/A _6999_/B _6563_/B _6479_/A vssd1 vssd1 vccd1 vccd1 _6575_/C sky130_fd_sc_hd__a211o_1
X_6451_ _6446_/B _6448_/B _6444_/Y vssd1 vssd1 vccd1 vccd1 _6452_/C sky130_fd_sc_hd__a21oi_1
X_6382_ _6384_/B _6382_/B _6382_/C vssd1 vssd1 vccd1 vccd1 _6383_/A sky130_fd_sc_hd__and3b_1
X_5402_ _5406_/B vssd1 vssd1 vccd1 vccd1 _5860_/A sky130_fd_sc_hd__clkbuf_2
X_8121_ _8233_/B _8121_/B vssd1 vssd1 vccd1 vccd1 _8125_/A sky130_fd_sc_hd__nor2_1
X_5333_ _5333_/A vssd1 vssd1 vccd1 vccd1 _5333_/X sky130_fd_sc_hd__clkbuf_2
X_5264_ _5294_/A vssd1 vssd1 vccd1 vccd1 _5264_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_8052_ _8052_/A _8052_/B vssd1 vssd1 vccd1 vccd1 _8053_/C sky130_fd_sc_hd__nand2_1
X_5195_ _8476_/Q _5205_/B vssd1 vssd1 vccd1 vccd1 _5195_/X sky130_fd_sc_hd__or2_1
X_7003_ _6507_/A _7001_/B _7184_/B _7002_/A vssd1 vssd1 vccd1 vccd1 _7003_/X sky130_fd_sc_hd__a22o_1
XFILLER_18_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7905_ _8142_/A vssd1 vssd1 vccd1 vccd1 _8054_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_36_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7836_ _7836_/A _8015_/B vssd1 vssd1 vccd1 vccd1 _8184_/A sky130_fd_sc_hd__xnor2_1
X_4979_ _5019_/B _5022_/B vssd1 vssd1 vccd1 vccd1 _5089_/B sky130_fd_sc_hd__or2_1
X_7767_ _7645_/B _7647_/B _7766_/Y vssd1 vssd1 vccd1 vccd1 _7978_/B sky130_fd_sc_hd__a21o_2
X_6718_ _6721_/B _7172_/A vssd1 vssd1 vccd1 vccd1 _6718_/X sky130_fd_sc_hd__or2b_1
X_7698_ _7951_/A _7742_/A vssd1 vssd1 vccd1 vccd1 _7699_/B sky130_fd_sc_hd__nand2_1
X_6649_ _6522_/X _6649_/B vssd1 vssd1 vccd1 vccd1 _6682_/B sky130_fd_sc_hd__and2b_2
X_8319_ _8319_/A _8319_/B vssd1 vssd1 vccd1 vccd1 _8332_/A sky130_fd_sc_hd__xor2_1
XFILLER_78_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8635__51 vssd1 vssd1 vccd1 vccd1 _8635__51/HI _8744_/A sky130_fd_sc_hd__conb_1
XFILLER_65_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5951_ _5951_/A _6153_/B vssd1 vssd1 vccd1 vccd1 _6037_/B sky130_fd_sc_hd__xnor2_1
XFILLER_37_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4902_ _4913_/A _5028_/D vssd1 vssd1 vccd1 vccd1 _5071_/C sky130_fd_sc_hd__or2_1
XFILLER_52_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5882_ _5880_/Y _5882_/B vssd1 vssd1 vccd1 vccd1 _5914_/B sky130_fd_sc_hd__and2b_1
X_4833_ _4592_/A _4830_/Y _4935_/A vssd1 vssd1 vccd1 vccd1 _4833_/X sky130_fd_sc_hd__o21a_1
X_7621_ _7621_/A _7621_/B vssd1 vssd1 vccd1 vccd1 _7744_/B sky130_fd_sc_hd__xnor2_1
XFILLER_33_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4764_ _4740_/C _4742_/B _4737_/A vssd1 vssd1 vccd1 vccd1 _4765_/B sky130_fd_sc_hd__a21oi_1
XFILLER_21_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7552_ _7616_/A _7552_/B vssd1 vssd1 vccd1 vccd1 _7562_/A sky130_fd_sc_hd__and2_1
X_6503_ _6584_/A _6632_/A vssd1 vssd1 vccd1 vccd1 _6585_/C sky130_fd_sc_hd__or2_1
X_7483_ _7483_/A _7487_/B vssd1 vssd1 vccd1 vccd1 _7484_/B sky130_fd_sc_hd__nand2_1
X_6434_ _6435_/A _6435_/B vssd1 vssd1 vccd1 vccd1 _6434_/Y sky130_fd_sc_hd__nor2_1
X_4695_ _5370_/A _4695_/B _4695_/C vssd1 vssd1 vccd1 vccd1 _4696_/A sky130_fd_sc_hd__and3_1
X_6365_ _6365_/A vssd1 vssd1 vccd1 vccd1 _8538_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8104_ _8104_/A _8224_/A vssd1 vssd1 vccd1 vccd1 _8108_/A sky130_fd_sc_hd__xnor2_1
X_6296_ _5333_/X _6295_/Y _6293_/A _4511_/B vssd1 vssd1 vccd1 vccd1 _8525_/D sky130_fd_sc_hd__o2bb2a_1
X_5316_ _8511_/Q vssd1 vssd1 vccd1 vccd1 _5339_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_5247_ _8489_/Q _6396_/B _5240_/B _8491_/Q vssd1 vssd1 vccd1 vccd1 _5248_/B sky130_fd_sc_hd__a31o_1
X_8035_ _8115_/A _8035_/B vssd1 vssd1 vccd1 vccd1 _8086_/B sky130_fd_sc_hd__and2_1
X_5178_ _5180_/B _5178_/B vssd1 vssd1 vccd1 vccd1 _5178_/Y sky130_fd_sc_hd__nand2_1
XFILLER_28_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7819_ _7781_/A _7781_/B _7818_/X vssd1 vssd1 vccd1 vccd1 _7872_/B sky130_fd_sc_hd__o21ai_1
XFILLER_12_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4480_ _8482_/Q _4480_/B vssd1 vssd1 vccd1 vccd1 _4481_/A sky130_fd_sc_hd__and2_1
XFILLER_7_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6150_ _6150_/A vssd1 vssd1 vccd1 vccd1 _6150_/Y sky130_fd_sc_hd__inv_2
X_5101_ _5085_/X _5088_/C _5101_/S vssd1 vssd1 vccd1 vccd1 _5102_/D sky130_fd_sc_hd__mux2_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6081_ _6081_/A _6081_/B vssd1 vssd1 vccd1 vccd1 _6232_/A sky130_fd_sc_hd__nor2_1
X_5032_ _5109_/C _5030_/X _5031_/X _4842_/C vssd1 vssd1 vccd1 vccd1 _5033_/D sky130_fd_sc_hd__o22a_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6983_ _6983_/A _6983_/B vssd1 vssd1 vccd1 vccd1 _6985_/B sky130_fd_sc_hd__xnor2_1
XFILLER_53_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8722_ _8722_/A _4306_/Y vssd1 vssd1 vccd1 vccd1 io_out[7] sky130_fd_sc_hd__ebufn_8
X_5934_ _5935_/A _5935_/B vssd1 vssd1 vccd1 vccd1 _6008_/A sky130_fd_sc_hd__nand2_1
X_5865_ _5866_/A _6129_/A vssd1 vssd1 vccd1 vccd1 _5924_/A sky130_fd_sc_hd__nand2_2
X_4816_ _5090_/A _5031_/C vssd1 vssd1 vccd1 vccd1 _5171_/C sky130_fd_sc_hd__or2_1
XFILLER_21_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7604_ _7604_/A _7604_/B vssd1 vssd1 vccd1 vccd1 _7725_/C sky130_fd_sc_hd__xor2_4
XFILLER_21_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5796_ _5528_/B _5530_/B _5564_/B _5646_/Y vssd1 vssd1 vccd1 vccd1 _5978_/B sky130_fd_sc_hd__a211o_1
X_8584_ input3/X _8584_/D vssd1 vssd1 vccd1 vccd1 _8584_/Q sky130_fd_sc_hd__dfxtp_1
X_4747_ _4747_/A _4798_/B vssd1 vssd1 vccd1 vccd1 _4996_/A sky130_fd_sc_hd__nor2_2
X_7535_ _7695_/B vssd1 vssd1 vccd1 vccd1 _8023_/A sky130_fd_sc_hd__clkbuf_2
X_4678_ _4684_/A vssd1 vssd1 vccd1 vccd1 _5207_/A sky130_fd_sc_hd__buf_2
X_7466_ _8573_/Q _7481_/B vssd1 vssd1 vccd1 vccd1 _7466_/X sky130_fd_sc_hd__xor2_1
X_6417_ _8552_/Q vssd1 vssd1 vccd1 vccd1 _6439_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7397_ _7398_/A _7398_/B vssd1 vssd1 vccd1 vccd1 _7409_/S sky130_fd_sc_hd__or2_1
X_6348_ _6389_/B vssd1 vssd1 vccd1 vccd1 _6348_/X sky130_fd_sc_hd__buf_2
XFILLER_88_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6279_ _6274_/B _5332_/X _5333_/A _6278_/Y vssd1 vssd1 vccd1 vccd1 _8522_/D sky130_fd_sc_hd__a22o_1
XFILLER_88_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8018_ _8012_/A _8012_/B _8011_/A vssd1 vssd1 vccd1 vccd1 _8082_/A sky130_fd_sc_hd__o21ai_1
XFILLER_56_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8605__21 vssd1 vssd1 vccd1 vccd1 _8605__21/HI _8700_/A sky130_fd_sc_hd__conb_1
XFILLER_94_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5650_ _5650_/A vssd1 vssd1 vccd1 vccd1 _5800_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4601_ _4645_/B vssd1 vssd1 vccd1 vccd1 _4657_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_5581_ _5581_/A _5581_/B vssd1 vssd1 vccd1 vccd1 _6243_/A sky130_fd_sc_hd__nand2_1
XFILLER_30_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7320_ _6873_/A _6873_/B _7319_/X vssd1 vssd1 vccd1 vccd1 _7331_/A sky130_fd_sc_hd__o21ai_1
XFILLER_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4532_ _4532_/A _4532_/B vssd1 vssd1 vccd1 vccd1 _8438_/D sky130_fd_sc_hd__nor2_1
X_7251_ _6509_/A _6509_/B _6505_/A _6505_/B vssd1 vssd1 vccd1 vccd1 _7358_/B sky130_fd_sc_hd__o2bb2a_1
X_4463_ _4735_/A _4759_/A _4882_/A _4748_/D vssd1 vssd1 vccd1 vccd1 _4805_/A sky130_fd_sc_hd__or4b_4
X_6202_ _5499_/A _5499_/C _5496_/B vssd1 vssd1 vccd1 vccd1 _6204_/A sky130_fd_sc_hd__a21oi_2
X_7182_ _7205_/A _7182_/B vssd1 vssd1 vccd1 vccd1 _7186_/A sky130_fd_sc_hd__xnor2_2
X_4394_ _5441_/B vssd1 vssd1 vccd1 vccd1 _4949_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6133_ _6131_/X _6133_/B vssd1 vssd1 vccd1 vccd1 _6134_/B sky130_fd_sc_hd__and2b_1
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6064_ _6075_/A _6075_/B _6076_/B vssd1 vssd1 vccd1 vccd1 _6078_/B sky130_fd_sc_hd__and3_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5015_ _5092_/D _5012_/X _5014_/X _4989_/A vssd1 vssd1 vccd1 vccd1 _5015_/X sky130_fd_sc_hd__o22a_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6966_ _7176_/A _7032_/B vssd1 vssd1 vccd1 vccd1 _7034_/S sky130_fd_sc_hd__nor2_2
XFILLER_53_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8705_ _8705_/A _4286_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[22] sky130_fd_sc_hd__ebufn_8
X_5917_ _5872_/A _5872_/B _5916_/X vssd1 vssd1 vccd1 vccd1 _5967_/A sky130_fd_sc_hd__a21boi_1
X_6897_ _6897_/A _6897_/B vssd1 vssd1 vccd1 vccd1 _6899_/B sky130_fd_sc_hd__xor2_2
XFILLER_21_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5848_ _6141_/A vssd1 vssd1 vccd1 vccd1 _5851_/A sky130_fd_sc_hd__inv_2
X_8567_ input3/X _8567_/D vssd1 vssd1 vccd1 vccd1 _8567_/Q sky130_fd_sc_hd__dfxtp_1
X_5779_ _5734_/A _5733_/B _5778_/X vssd1 vssd1 vccd1 vccd1 _5780_/B sky130_fd_sc_hd__o21ai_4
XFILLER_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7518_ _7518_/A _7518_/B vssd1 vssd1 vccd1 vccd1 _7542_/A sky130_fd_sc_hd__or2_1
X_8498_ input3/X _8498_/D vssd1 vssd1 vccd1 vccd1 _8498_/Q sky130_fd_sc_hd__dfxtp_1
X_7449_ _7494_/A _7448_/X _6462_/A vssd1 vssd1 vccd1 vccd1 _7449_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_88_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6820_ _6721_/A _7122_/C _6679_/B vssd1 vssd1 vccd1 vccd1 _7286_/B sky130_fd_sc_hd__o21ai_2
XFILLER_90_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6751_ _6751_/A _6751_/B vssd1 vssd1 vccd1 vccd1 _7032_/A sky130_fd_sc_hd__or2_1
X_6682_ _6682_/A _6682_/B vssd1 vssd1 vccd1 vccd1 _7001_/B sky130_fd_sc_hd__xor2_4
X_5702_ _6053_/A _6053_/B vssd1 vssd1 vccd1 vccd1 _5715_/A sky130_fd_sc_hd__and2_1
X_5633_ _5633_/A _5633_/B _5632_/X vssd1 vssd1 vccd1 vccd1 _5720_/B sky130_fd_sc_hd__or3b_1
X_8421_ _8421_/A _8429_/S vssd1 vssd1 vccd1 vccd1 _8425_/A sky130_fd_sc_hd__or2b_1
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8352_ _8352_/A _8352_/B vssd1 vssd1 vccd1 vccd1 _8353_/B sky130_fd_sc_hd__xnor2_4
X_5564_ _5978_/A _5564_/B vssd1 vssd1 vccd1 vccd1 _5980_/C sky130_fd_sc_hd__nand2_1
X_7303_ _7303_/A _7303_/B vssd1 vssd1 vccd1 vccd1 _7309_/A sky130_fd_sc_hd__xnor2_1
X_4515_ _8434_/Q _8433_/Q vssd1 vssd1 vccd1 vccd1 _4516_/C sky130_fd_sc_hd__nand2_1
X_8283_ _8163_/A _8163_/B _8282_/X vssd1 vssd1 vccd1 vccd1 _8339_/A sky130_fd_sc_hd__o21a_1
X_5495_ _5495_/A _8463_/Q vssd1 vssd1 vccd1 vccd1 _5496_/B sky130_fd_sc_hd__or2_1
X_7234_ _7234_/A _7234_/B vssd1 vssd1 vccd1 vccd1 _7236_/B sky130_fd_sc_hd__xnor2_1
X_4446_ _8457_/Q vssd1 vssd1 vccd1 vccd1 _6482_/B sky130_fd_sc_hd__buf_4
X_7165_ _7165_/A _7165_/B vssd1 vssd1 vccd1 vccd1 _7166_/B sky130_fd_sc_hd__xnor2_1
X_4377_ _4381_/A vssd1 vssd1 vccd1 vccd1 _4377_/Y sky130_fd_sc_hd__inv_2
X_6116_ _5987_/A _5987_/B _6115_/X vssd1 vssd1 vccd1 vccd1 _6117_/B sky130_fd_sc_hd__a21oi_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7096_ _7098_/B _7264_/A _7098_/A vssd1 vssd1 vccd1 vccd1 _7097_/B sky130_fd_sc_hd__o21ai_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6047_ _6095_/B _6047_/B vssd1 vssd1 vccd1 vccd1 _6048_/B sky130_fd_sc_hd__xnor2_1
XFILLER_37_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8596__12 vssd1 vssd1 vccd1 vccd1 _8596__12/HI _8691_/A sky130_fd_sc_hd__conb_1
XFILLER_81_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7998_ _8041_/A _7924_/B vssd1 vssd1 vccd1 vccd1 _7998_/X sky130_fd_sc_hd__or2b_1
X_6949_ _6949_/A _6949_/B vssd1 vssd1 vccd1 vccd1 _6949_/Y sky130_fd_sc_hd__nand2_1
XFILLER_53_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4300_ _4301_/A vssd1 vssd1 vccd1 vccd1 _4300_/Y sky130_fd_sc_hd__inv_2
X_5280_ _8501_/Q _5283_/C vssd1 vssd1 vccd1 vccd1 _5282_/A sky130_fd_sc_hd__and2_1
XFILLER_4_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8680__96 vssd1 vssd1 vccd1 vccd1 _8680__96/HI _8789_/A sky130_fd_sc_hd__conb_1
X_7921_ _7921_/A _7921_/B vssd1 vssd1 vccd1 vccd1 _8025_/A sky130_fd_sc_hd__nand2_1
XFILLER_82_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7852_ _7899_/A _8260_/B vssd1 vssd1 vccd1 vccd1 _8069_/A sky130_fd_sc_hd__nor2_1
XFILLER_90_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4995_ _5031_/B _5169_/B _4995_/C _5148_/C vssd1 vssd1 vccd1 vccd1 _4996_/C sky130_fd_sc_hd__or4_1
X_6803_ _6863_/B _6863_/C _6863_/A vssd1 vssd1 vccd1 vccd1 _6814_/A sky130_fd_sc_hd__a21bo_1
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7783_ _7783_/A _7783_/B vssd1 vssd1 vccd1 vccd1 _7783_/X sky130_fd_sc_hd__and2_1
X_6734_ _6804_/A _6616_/B _6616_/C vssd1 vssd1 vccd1 vccd1 _6740_/A sky130_fd_sc_hd__a21bo_1
XFILLER_51_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6665_ _6939_/A _6680_/A vssd1 vssd1 vccd1 vccd1 _6926_/A sky130_fd_sc_hd__nor2_1
X_8404_ _8404_/A vssd1 vssd1 vccd1 vccd1 _8583_/D sky130_fd_sc_hd__clkbuf_1
X_6596_ _6604_/A _6596_/B vssd1 vssd1 vccd1 vccd1 _6597_/B sky130_fd_sc_hd__nand2_1
X_5616_ _5499_/A _5496_/B _5499_/C _5494_/X vssd1 vssd1 vccd1 vccd1 _5767_/B sky130_fd_sc_hd__a31o_2
X_8335_ _8281_/A _8281_/B _8334_/Y vssd1 vssd1 vccd1 vccd1 _8336_/B sky130_fd_sc_hd__o21ai_1
X_5547_ _5547_/A _5547_/B vssd1 vssd1 vccd1 vccd1 _5548_/B sky130_fd_sc_hd__or2_1
X_8266_ _8266_/A _8266_/B vssd1 vssd1 vccd1 vccd1 _8267_/B sky130_fd_sc_hd__or2_1
XFILLER_2_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5478_ _6188_/A _5637_/A _5829_/C _5831_/A vssd1 vssd1 vccd1 vccd1 _5601_/B sky130_fd_sc_hd__o31ai_1
X_7217_ _7259_/A _7259_/B vssd1 vssd1 vccd1 vccd1 _7217_/Y sky130_fd_sc_hd__nand2_1
X_4429_ _4725_/A vssd1 vssd1 vccd1 vccd1 _4748_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8197_ _8207_/A _8207_/B _8196_/X vssd1 vssd1 vccd1 vccd1 _8211_/A sky130_fd_sc_hd__o21a_1
XFILLER_86_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7148_ _7152_/A _7148_/B vssd1 vssd1 vccd1 vccd1 _7181_/A sky130_fd_sc_hd__xor2_2
X_7079_ _7079_/A _7079_/B vssd1 vssd1 vccd1 vccd1 _7085_/B sky130_fd_sc_hd__xnor2_1
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4780_ _4780_/A _4780_/B _4899_/A vssd1 vssd1 vccd1 vccd1 _4994_/B sky130_fd_sc_hd__or3_2
X_6450_ _6455_/A _6450_/B vssd1 vssd1 vccd1 vccd1 _6459_/A sky130_fd_sc_hd__nand2_1
X_6381_ _8542_/Q _6380_/B _6375_/B _8544_/Q vssd1 vssd1 vccd1 vccd1 _6382_/C sky130_fd_sc_hd__a31o_1
X_5401_ _5855_/A vssd1 vssd1 vccd1 vccd1 _5406_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_8120_ _8120_/A _8120_/B vssd1 vssd1 vccd1 vccd1 _8121_/B sky130_fd_sc_hd__nor2_1
X_5332_ _5332_/A vssd1 vssd1 vccd1 vccd1 _5332_/X sky130_fd_sc_hd__clkbuf_2
X_5263_ _8496_/Q _5263_/B vssd1 vssd1 vccd1 vccd1 _5270_/C sky130_fd_sc_hd__and2_1
X_8051_ _7966_/A _7966_/B _8050_/X vssd1 vssd1 vccd1 vccd1 _8057_/A sky130_fd_sc_hd__a21bo_1
X_5194_ _5207_/A vssd1 vssd1 vccd1 vccd1 _5205_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_7002_ _7002_/A _7248_/B vssd1 vssd1 vccd1 vccd1 _7250_/A sky130_fd_sc_hd__nand2_2
XFILLER_68_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7904_ _7904_/A _7904_/B vssd1 vssd1 vccd1 vccd1 _7909_/A sky130_fd_sc_hd__xor2_4
XFILLER_24_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7835_ _8012_/A _7835_/B vssd1 vssd1 vccd1 vccd1 _8015_/B sky130_fd_sc_hd__nand2_1
XFILLER_51_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4978_ _5016_/A _5171_/A vssd1 vssd1 vccd1 vccd1 _5022_/C sky130_fd_sc_hd__or2_1
XFILLER_11_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7766_ _7766_/A _7766_/B vssd1 vssd1 vccd1 vccd1 _7766_/Y sky130_fd_sc_hd__nor2_1
X_6717_ _6721_/B _7172_/A vssd1 vssd1 vccd1 vccd1 _6938_/B sky130_fd_sc_hd__xor2_1
X_7697_ _7697_/A _7697_/B vssd1 vssd1 vccd1 vccd1 _8366_/A sky130_fd_sc_hd__nand2_1
X_6648_ _6574_/B _6575_/B _6575_/C _6521_/X vssd1 vssd1 vccd1 vccd1 _6682_/A sky130_fd_sc_hd__a31o_2
XFILLER_50_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6579_ _6939_/B _7323_/B _6786_/B vssd1 vssd1 vccd1 vccd1 _6580_/B sky130_fd_sc_hd__or3_2
X_8318_ _7961_/A _7734_/A _8053_/B _8317_/Y vssd1 vssd1 vccd1 vccd1 _8319_/B sky130_fd_sc_hd__o211a_1
X_8249_ _8249_/A _8249_/B vssd1 vssd1 vccd1 vccd1 _8306_/B sky130_fd_sc_hd__and2_1
XFILLER_47_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8650__66 vssd1 vssd1 vccd1 vccd1 _8650__66/HI _8759_/A sky130_fd_sc_hd__conb_1
XFILLER_92_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5950_ _6137_/A _5930_/A _6137_/B vssd1 vssd1 vccd1 vccd1 _6153_/B sky130_fd_sc_hd__a21o_1
X_4901_ _5107_/C _5055_/A _4915_/A vssd1 vssd1 vccd1 vccd1 _5028_/D sky130_fd_sc_hd__or3_1
XFILLER_52_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5881_ _5880_/A _5880_/C _5880_/B vssd1 vssd1 vccd1 vccd1 _5882_/B sky130_fd_sc_hd__o21ai_1
X_7620_ _7620_/A _7740_/A _7741_/A vssd1 vssd1 vccd1 vccd1 _7621_/B sky130_fd_sc_hd__or3_2
X_4832_ _5136_/A vssd1 vssd1 vccd1 vccd1 _4935_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_21_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4763_ _4779_/A _4791_/A _4908_/B _4811_/A vssd1 vssd1 vccd1 vccd1 _4886_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_21_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7551_ _8461_/Q _8585_/Q vssd1 vssd1 vccd1 vccd1 _7552_/B sky130_fd_sc_hd__or2b_1
X_6502_ _6534_/A _6751_/B vssd1 vssd1 vccd1 vccd1 _6632_/A sky130_fd_sc_hd__xnor2_2
X_4694_ _4698_/B _4698_/C vssd1 vssd1 vccd1 vccd1 _4695_/C sky130_fd_sc_hd__nand2_1
X_7482_ _7539_/A _7482_/B vssd1 vssd1 vccd1 vccd1 _7487_/B sky130_fd_sc_hd__or2_1
X_6433_ _6433_/A _8549_/Q vssd1 vssd1 vccd1 vccd1 _6435_/B sky130_fd_sc_hd__xor2_1
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6364_ _6366_/B _6364_/B _6382_/B vssd1 vssd1 vccd1 vccd1 _6365_/A sky130_fd_sc_hd__and3b_1
X_5315_ _8512_/Q vssd1 vssd1 vccd1 vccd1 _5345_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_8103_ _8227_/A _8225_/B vssd1 vssd1 vccd1 vccd1 _8224_/A sky130_fd_sc_hd__xor2_1
X_6295_ _6295_/A _6295_/B vssd1 vssd1 vccd1 vccd1 _6295_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_88_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5246_ _8491_/Q _8490_/Q _5246_/C vssd1 vssd1 vccd1 vccd1 _5253_/C sky130_fd_sc_hd__and3_1
X_8034_ _8034_/A _8034_/B vssd1 vssd1 vccd1 vccd1 _8035_/B sky130_fd_sc_hd__or2_1
XFILLER_29_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5177_ _4790_/B _4800_/A _4765_/A _4466_/B _4755_/A vssd1 vssd1 vccd1 vccd1 _5185_/A
+ sky130_fd_sc_hd__a2111o_1
XFILLER_83_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7818_ _7818_/A _7818_/B vssd1 vssd1 vccd1 vccd1 _7818_/X sky130_fd_sc_hd__or2_1
X_7749_ _7750_/A _7750_/B _7750_/C vssd1 vssd1 vccd1 vccd1 _7838_/A sky130_fd_sc_hd__a21o_1
XFILLER_10_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5100_ _4873_/A _5107_/C _5053_/B _5033_/C _5099_/X vssd1 vssd1 vccd1 vccd1 _5100_/X
+ sky130_fd_sc_hd__o32a_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6080_ _6079_/A _6079_/C _6079_/B vssd1 vssd1 vccd1 vccd1 _6081_/B sky130_fd_sc_hd__o21a_1
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5031_ _5093_/A _5031_/B _5031_/C _5136_/C vssd1 vssd1 vccd1 vccd1 _5031_/X sky130_fd_sc_hd__or4_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8721_ _8721_/A _4305_/Y vssd1 vssd1 vccd1 vccd1 io_out[6] sky130_fd_sc_hd__ebufn_8
X_6982_ _7050_/A _7050_/B vssd1 vssd1 vccd1 vccd1 _6985_/A sky130_fd_sc_hd__nand2_1
XFILLER_80_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5933_ _5846_/Y _6200_/A _6125_/A vssd1 vssd1 vccd1 vccd1 _5935_/B sky130_fd_sc_hd__o21ba_1
X_5864_ _5918_/A _5992_/A _5918_/C vssd1 vssd1 vccd1 vccd1 _6129_/A sky130_fd_sc_hd__nand3_2
XFILLER_33_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4815_ _4969_/B _4886_/D vssd1 vssd1 vccd1 vccd1 _5031_/C sky130_fd_sc_hd__or2_1
X_7603_ _7552_/B _7576_/A _7562_/C _7602_/Y vssd1 vssd1 vccd1 vccd1 _7604_/B sky130_fd_sc_hd__a31o_1
X_8583_ input3/X _8583_/D vssd1 vssd1 vccd1 vccd1 _8583_/Q sky130_fd_sc_hd__dfxtp_1
X_5795_ _5795_/A vssd1 vssd1 vccd1 vccd1 _5918_/A sky130_fd_sc_hd__clkbuf_2
X_7534_ _7679_/A _7532_/B _7533_/X vssd1 vssd1 vccd1 vccd1 _7549_/A sky130_fd_sc_hd__a21bo_1
X_4746_ _4796_/B vssd1 vssd1 vccd1 vccd1 _4798_/B sky130_fd_sc_hd__buf_2
X_4677_ _4670_/A _4735_/B _4882_/A _4780_/A vssd1 vssd1 vccd1 vccd1 _4677_/X sky130_fd_sc_hd__a31o_1
X_7465_ _7465_/A vssd1 vssd1 vccd1 vccd1 _8572_/D sky130_fd_sc_hd__clkbuf_1
X_7396_ _7391_/B _7393_/B _7391_/A vssd1 vssd1 vccd1 vccd1 _7398_/B sky130_fd_sc_hd__a21bo_1
X_6416_ _6445_/B vssd1 vssd1 vccd1 vccd1 _6450_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6347_ _6351_/A _6351_/C vssd1 vssd1 vccd1 vccd1 _6350_/A sky130_fd_sc_hd__and2_1
XFILLER_88_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6278_ _6278_/A _6278_/B vssd1 vssd1 vccd1 vccd1 _6278_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_69_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5229_ _5260_/A vssd1 vssd1 vccd1 vccd1 _5230_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_29_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8017_ _8188_/A _8188_/B vssd1 vssd1 vccd1 vccd1 _8190_/B sky130_fd_sc_hd__nor2_1
XFILLER_84_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8620__36 vssd1 vssd1 vccd1 vccd1 _8620__36/HI _8715_/A sky130_fd_sc_hd__conb_1
XFILLER_35_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4600_ _6427_/A _4671_/B vssd1 vssd1 vccd1 vccd1 _4645_/B sky130_fd_sc_hd__nor2_1
X_5580_ _5978_/A _6244_/B _5705_/A vssd1 vssd1 vccd1 vccd1 _5581_/B sky130_fd_sc_hd__a21oi_1
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4531_ _8438_/Q _4533_/C _4524_/X vssd1 vssd1 vccd1 vccd1 _4532_/B sky130_fd_sc_hd__o21ai_1
X_7250_ _7250_/A _7250_/B vssd1 vssd1 vccd1 vccd1 _7358_/A sky130_fd_sc_hd__xor2_1
X_4462_ _4759_/B vssd1 vssd1 vccd1 vccd1 _4882_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6201_ _6201_/A _6201_/B vssd1 vssd1 vccd1 vccd1 _6208_/A sky130_fd_sc_hd__xnor2_1
X_7181_ _7181_/A _7181_/B vssd1 vssd1 vccd1 vccd1 _7182_/B sky130_fd_sc_hd__xnor2_2
X_4393_ _8458_/Q vssd1 vssd1 vccd1 vccd1 _5441_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_58_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6132_ _6132_/A _6132_/B _6132_/C vssd1 vssd1 vccd1 vccd1 _6133_/B sky130_fd_sc_hd__or3_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6063_ _6063_/A _6063_/B vssd1 vssd1 vccd1 vccd1 _6076_/B sky130_fd_sc_hd__xnor2_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5014_ _5160_/C _5064_/C _5033_/C _5014_/D vssd1 vssd1 vccd1 vccd1 _5014_/X sky130_fd_sc_hd__or4_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6965_ _6972_/A _6964_/B _6736_/B _6751_/A vssd1 vssd1 vccd1 vccd1 _7044_/B sky130_fd_sc_hd__o22ai_4
X_8704_ _8704_/A _4285_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[21] sky130_fd_sc_hd__ebufn_8
XFILLER_53_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5916_ _5916_/A _5854_/B vssd1 vssd1 vccd1 vccd1 _5916_/X sky130_fd_sc_hd__or2b_1
X_6896_ _6896_/A _6896_/B _6896_/C vssd1 vssd1 vccd1 vccd1 _6899_/A sky130_fd_sc_hd__nand3_1
XFILLER_34_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5847_ _6021_/A _5767_/X _5846_/Y vssd1 vssd1 vccd1 vccd1 _6141_/A sky130_fd_sc_hd__a21o_1
X_8566_ input3/X _8566_/D vssd1 vssd1 vccd1 vccd1 _8566_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5778_ _5778_/A _5942_/B vssd1 vssd1 vccd1 vccd1 _5778_/X sky130_fd_sc_hd__or2_2
X_4729_ _4790_/A _4790_/B _4773_/A vssd1 vssd1 vccd1 vccd1 _5153_/B sky130_fd_sc_hd__nor3_2
X_8497_ input3/X _8497_/D vssd1 vssd1 vccd1 vccd1 _8497_/Q sky130_fd_sc_hd__dfxtp_1
X_7517_ _7518_/A _7518_/B vssd1 vssd1 vccd1 vccd1 _7517_/X sky130_fd_sc_hd__and2_1
X_7448_ _8430_/A vssd1 vssd1 vccd1 vccd1 _7448_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_89_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7379_ _8548_/Q _7380_/A vssd1 vssd1 vccd1 vccd1 _7381_/A sky130_fd_sc_hd__or2b_1
XFILLER_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6750_ _6980_/A _7291_/B _6749_/Y vssd1 vssd1 vccd1 vccd1 _6875_/B sky130_fd_sc_hd__a21bo_1
XFILLER_35_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5701_ _5812_/B _5747_/B _5748_/B vssd1 vssd1 vccd1 vccd1 _5717_/A sky130_fd_sc_hd__and3_1
X_6681_ _7323_/A _6784_/A vssd1 vssd1 vccd1 vccd1 _6688_/A sky130_fd_sc_hd__or2_1
X_8420_ _8420_/A vssd1 vssd1 vccd1 vccd1 _8585_/D sky130_fd_sc_hd__clkbuf_1
X_5632_ _5719_/A _5632_/B vssd1 vssd1 vccd1 vccd1 _5632_/X sky130_fd_sc_hd__and2_1
X_8351_ _8351_/A _8351_/B vssd1 vssd1 vccd1 vccd1 _8352_/B sky130_fd_sc_hd__xnor2_2
X_5563_ _5563_/A _5563_/B vssd1 vssd1 vccd1 vccd1 _5564_/B sky130_fd_sc_hd__xor2_1
X_4514_ _4536_/A vssd1 vssd1 vccd1 vccd1 _4575_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7302_ _7302_/A _7302_/B vssd1 vssd1 vccd1 vccd1 _7303_/B sky130_fd_sc_hd__xnor2_1
X_8282_ _8282_/A _8282_/B vssd1 vssd1 vccd1 vccd1 _8282_/X sky130_fd_sc_hd__or2_1
X_5494_ _5495_/A _7613_/B vssd1 vssd1 vccd1 vccd1 _5494_/X sky130_fd_sc_hd__and2_1
X_4445_ _4445_/A vssd1 vssd1 vccd1 vccd1 _8727_/A sky130_fd_sc_hd__clkbuf_1
X_7233_ _7233_/A _7233_/B _7233_/C vssd1 vssd1 vccd1 vccd1 _7247_/A sky130_fd_sc_hd__or3_1
X_4376_ _4382_/A vssd1 vssd1 vccd1 vccd1 _4381_/A sky130_fd_sc_hd__clkbuf_2
X_7164_ _7193_/A _7193_/B _7194_/B _7163_/X vssd1 vssd1 vccd1 vccd1 _7167_/A sky130_fd_sc_hd__a31oi_2
X_6115_ _5988_/B _6115_/B vssd1 vssd1 vccd1 vccd1 _6115_/X sky130_fd_sc_hd__and2b_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7095_ _7272_/C _7095_/B vssd1 vssd1 vccd1 vccd1 _7098_/A sky130_fd_sc_hd__and2_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6046_ _6046_/A _6046_/B vssd1 vssd1 vccd1 vccd1 _6047_/B sky130_fd_sc_hd__xnor2_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7997_ _7933_/A _7933_/B _7934_/A vssd1 vssd1 vccd1 vccd1 _8010_/A sky130_fd_sc_hd__a21oi_1
X_6948_ _6948_/A _7015_/A vssd1 vssd1 vccd1 vccd1 _6953_/A sky130_fd_sc_hd__or2b_1
X_6879_ _6879_/A _6879_/B _6879_/C vssd1 vssd1 vccd1 vccd1 _6883_/A sky130_fd_sc_hd__nand3_1
XFILLER_10_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8549_ input3/X _8549_/D vssd1 vssd1 vccd1 vccd1 _8549_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7920_ _8231_/A vssd1 vssd1 vccd1 vccd1 _8041_/C sky130_fd_sc_hd__clkbuf_2
X_7851_ _8147_/B vssd1 vssd1 vccd1 vccd1 _8260_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6802_ _6980_/B _6802_/B _6802_/C vssd1 vssd1 vccd1 vccd1 _6863_/A sky130_fd_sc_hd__nand3_1
X_4994_ _5104_/A _4994_/B vssd1 vssd1 vccd1 vccd1 _5148_/C sky130_fd_sc_hd__nand2_2
X_7782_ _7783_/A _7783_/B vssd1 vssd1 vccd1 vccd1 _7782_/Y sky130_fd_sc_hd__nor2_1
X_6733_ _6733_/A _6733_/B vssd1 vssd1 vccd1 vccd1 _6879_/B sky130_fd_sc_hd__nand2_1
X_6664_ _6930_/A _6902_/B _6663_/Y vssd1 vssd1 vccd1 vccd1 _6731_/A sky130_fd_sc_hd__o21a_1
X_5615_ _5615_/A _5724_/A vssd1 vssd1 vccd1 vccd1 _5618_/A sky130_fd_sc_hd__nor2_1
X_8403_ _8403_/A _8403_/B vssd1 vssd1 vccd1 vccd1 _8404_/A sky130_fd_sc_hd__and2_1
X_6595_ _6595_/A _6543_/X vssd1 vssd1 vccd1 vccd1 _6597_/A sky130_fd_sc_hd__or2b_1
XFILLER_3_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8334_ _8334_/A _8334_/B vssd1 vssd1 vccd1 vccd1 _8334_/Y sky130_fd_sc_hd__nand2_1
X_5546_ _5547_/A _5547_/B vssd1 vssd1 vccd1 vccd1 _5548_/A sky130_fd_sc_hd__nand2_1
X_8265_ _8266_/A _8266_/B vssd1 vssd1 vccd1 vccd1 _8267_/A sky130_fd_sc_hd__nand2_1
X_5477_ _6188_/B _5932_/A vssd1 vssd1 vccd1 vccd1 _5831_/A sky130_fd_sc_hd__or2_2
X_7216_ _7226_/A _7213_/B _7215_/X vssd1 vssd1 vccd1 vccd1 _7259_/B sky130_fd_sc_hd__a21oi_1
X_4428_ _7494_/B vssd1 vssd1 vccd1 vccd1 _4725_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_8656__72 vssd1 vssd1 vccd1 vccd1 _8656__72/HI _8765_/A sky130_fd_sc_hd__conb_1
X_8196_ _8196_/A _8196_/B vssd1 vssd1 vccd1 vccd1 _8196_/X sky130_fd_sc_hd__or2_1
X_7147_ _7146_/B _7146_/C _7146_/A vssd1 vssd1 vccd1 vccd1 _7345_/B sky130_fd_sc_hd__a21oi_1
XFILLER_86_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4359_ _4363_/A vssd1 vssd1 vccd1 vccd1 _4359_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7078_ _7109_/A _7109_/B _7060_/B _7077_/Y vssd1 vssd1 vccd1 vccd1 _7085_/A sky130_fd_sc_hd__a31o_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6029_ _5637_/B _5942_/B _5943_/B _5943_/A vssd1 vssd1 vccd1 vccd1 _6030_/B sky130_fd_sc_hd__o22a_1
XFILLER_73_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6380_ _8544_/Q _6380_/B _6380_/C vssd1 vssd1 vccd1 vccd1 _6384_/B sky130_fd_sc_hd__and3_1
X_5400_ _5400_/A _5400_/B vssd1 vssd1 vccd1 vccd1 _5855_/A sky130_fd_sc_hd__xnor2_4
X_5331_ _5331_/A vssd1 vssd1 vccd1 vccd1 _8509_/D sky130_fd_sc_hd__clkbuf_1
X_8050_ _8050_/A _7965_/B vssd1 vssd1 vccd1 vccd1 _8050_/X sky130_fd_sc_hd__or2b_1
XFILLER_87_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7001_ _7248_/A _7001_/B vssd1 vssd1 vccd1 vccd1 _7116_/B sky130_fd_sc_hd__nand2_2
X_5262_ _5262_/A vssd1 vssd1 vccd1 vccd1 _8495_/D sky130_fd_sc_hd__clkbuf_1
X_5193_ _8517_/Q _5188_/X _5192_/X _6426_/A vssd1 vssd1 vccd1 vccd1 _8475_/D sky130_fd_sc_hd__o211a_1
XFILLER_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7903_ _7903_/A _7903_/B vssd1 vssd1 vccd1 vccd1 _7904_/B sky130_fd_sc_hd__xor2_4
XFILLER_34_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7834_ _7834_/A _7834_/B vssd1 vssd1 vccd1 vccd1 _7835_/B sky130_fd_sc_hd__or2_1
XFILLER_36_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7765_ _7805_/A _7803_/A vssd1 vssd1 vccd1 vccd1 _7778_/A sky130_fd_sc_hd__nand2_1
X_4977_ _5146_/A _5074_/A _4977_/C _5009_/C vssd1 vssd1 vccd1 vccd1 _4977_/X sky130_fd_sc_hd__or4_1
X_6716_ _6647_/A _7116_/A _6987_/B _7054_/A vssd1 vssd1 vccd1 vccd1 _7172_/A sky130_fd_sc_hd__o22ai_4
XFILLER_51_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7696_ _8099_/A _8367_/B _7824_/A vssd1 vssd1 vccd1 vccd1 _7697_/B sky130_fd_sc_hd__a21oi_1
X_6647_ _6647_/A _6647_/B vssd1 vssd1 vccd1 vccd1 _6658_/A sky130_fd_sc_hd__xnor2_1
X_6578_ _7069_/B vssd1 vssd1 vccd1 vccd1 _6786_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_8317_ _8317_/A _8317_/B vssd1 vssd1 vccd1 vccd1 _8317_/Y sky130_fd_sc_hd__nand2_1
X_5529_ _5422_/A _5419_/Y _5422_/B _5420_/A vssd1 vssd1 vccd1 vccd1 _5530_/B sky130_fd_sc_hd__a31o_1
XFILLER_59_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8248_ _8248_/A _8248_/B vssd1 vssd1 vccd1 vccd1 _8255_/B sky130_fd_sc_hd__and2_1
XFILLER_78_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8179_ _7788_/B _7788_/C _7788_/A vssd1 vssd1 vccd1 vccd1 _8181_/A sky130_fd_sc_hd__a21boi_2
XFILLER_59_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4900_ _4991_/A _4906_/D _5041_/C vssd1 vssd1 vccd1 vccd1 _4900_/X sky130_fd_sc_hd__or3_1
XFILLER_80_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5880_ _5880_/A _5880_/B _5880_/C vssd1 vssd1 vccd1 vccd1 _5880_/Y sky130_fd_sc_hd__nor3_1
X_4831_ _5064_/A vssd1 vssd1 vccd1 vccd1 _5136_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_33_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4762_ _4762_/A _4766_/B _4762_/C vssd1 vssd1 vccd1 vccd1 _4811_/A sky130_fd_sc_hd__nor3_1
XFILLER_60_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7550_ _8585_/Q _6521_/B vssd1 vssd1 vccd1 vccd1 _7616_/A sky130_fd_sc_hd__or2b_1
X_6501_ _6501_/A _6501_/B vssd1 vssd1 vccd1 vccd1 _6751_/B sky130_fd_sc_hd__xnor2_2
X_4693_ _4698_/B _4698_/C vssd1 vssd1 vccd1 vccd1 _4695_/B sky130_fd_sc_hd__or2_1
X_7481_ _7539_/A _7481_/B vssd1 vssd1 vccd1 vccd1 _7483_/A sky130_fd_sc_hd__nand2_1
X_6432_ _6432_/A vssd1 vssd1 vccd1 vccd1 _6432_/X sky130_fd_sc_hd__clkbuf_2
X_6363_ _6362_/B _8536_/Q _6356_/A _8538_/Q vssd1 vssd1 vccd1 vccd1 _6364_/B sky130_fd_sc_hd__a31o_1
X_8102_ _8105_/B _8102_/B _8229_/B vssd1 vssd1 vccd1 vccd1 _8225_/B sky130_fd_sc_hd__and3b_1
X_6294_ _6294_/A _6297_/B vssd1 vssd1 vccd1 vccd1 _6295_/B sky130_fd_sc_hd__nor2_1
X_5314_ _8510_/Q vssd1 vssd1 vccd1 vccd1 _5335_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5245_ _6396_/B _5246_/C _5244_/Y vssd1 vssd1 vccd1 vccd1 _8490_/D sky130_fd_sc_hd__a21oi_1
X_8033_ _8034_/A _8034_/B vssd1 vssd1 vccd1 vccd1 _8115_/A sky130_fd_sc_hd__nand2_1
X_8626__42 vssd1 vssd1 vccd1 vccd1 _8626__42/HI _8721_/A sky130_fd_sc_hd__conb_1
XFILLER_29_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5176_ _5141_/X _5175_/X _5176_/S vssd1 vssd1 vccd1 vccd1 _5176_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7817_ _7817_/A _7817_/B vssd1 vssd1 vccd1 vccd1 _7871_/B sky130_fd_sc_hd__nand2_1
X_7748_ _7866_/A _7748_/B vssd1 vssd1 vccd1 vccd1 _7750_/C sky130_fd_sc_hd__nand2_1
X_7679_ _7679_/A _8023_/A vssd1 vssd1 vccd1 vccd1 _7694_/A sky130_fd_sc_hd__nand2_1
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5030_ _5104_/A _5030_/B _5030_/C _5041_/C vssd1 vssd1 vccd1 vccd1 _5030_/X sky130_fd_sc_hd__or4_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6981_ _7176_/A _6978_/A _6981_/S vssd1 vssd1 vccd1 vccd1 _7050_/B sky130_fd_sc_hd__mux2_1
X_8720_ _8720_/A _4304_/Y vssd1 vssd1 vccd1 vccd1 io_out[5] sky130_fd_sc_hd__ebufn_8
XFILLER_65_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5932_ _5932_/A _5932_/B vssd1 vssd1 vccd1 vccd1 _6125_/A sky130_fd_sc_hd__nor2_1
XFILLER_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5863_ _5863_/A _5863_/B vssd1 vssd1 vccd1 vccd1 _5866_/A sky130_fd_sc_hd__xor2_1
X_4814_ _4985_/A _4869_/B vssd1 vssd1 vccd1 vccd1 _4886_/D sky130_fd_sc_hd__or2_1
XFILLER_61_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5794_ _5794_/A _6226_/A vssd1 vssd1 vccd1 vccd1 _5809_/C sky130_fd_sc_hd__xnor2_1
X_7602_ _7616_/A vssd1 vssd1 vccd1 vccd1 _7602_/Y sky130_fd_sc_hd__inv_2
X_8582_ input3/X _8582_/D vssd1 vssd1 vccd1 vccd1 _8582_/Q sky130_fd_sc_hd__dfxtp_2
X_4745_ _5099_/C _5160_/C vssd1 vssd1 vccd1 vccd1 _4855_/A sky130_fd_sc_hd__or2_1
X_7533_ _7682_/A _7682_/B vssd1 vssd1 vccd1 vccd1 _7533_/X sky130_fd_sc_hd__or2_1
XFILLER_31_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4676_ _4676_/A vssd1 vssd1 vccd1 vccd1 _4808_/A sky130_fd_sc_hd__clkbuf_2
X_7464_ _8403_/A _7464_/B vssd1 vssd1 vccd1 vccd1 _7465_/A sky130_fd_sc_hd__and2_1
X_6415_ _8549_/Q vssd1 vssd1 vccd1 vccd1 _6445_/B sky130_fd_sc_hd__inv_2
X_7395_ _8565_/Q _7403_/B vssd1 vssd1 vccd1 vccd1 _7398_/A sky130_fd_sc_hd__xor2_1
X_6346_ _6346_/A vssd1 vssd1 vccd1 vccd1 _8532_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6277_ _6267_/S _6272_/B _6271_/A vssd1 vssd1 vccd1 vccd1 _6278_/B sky130_fd_sc_hd__o21a_1
X_8016_ _8016_/A _8016_/B vssd1 vssd1 vccd1 vccd1 _8188_/B sky130_fd_sc_hd__xnor2_1
X_5228_ _6328_/A _6465_/A vssd1 vssd1 vccd1 vccd1 _5260_/A sky130_fd_sc_hd__and2_1
X_5159_ _5162_/B _5159_/B vssd1 vssd1 vccd1 vccd1 _5159_/X sky130_fd_sc_hd__or2_1
XFILLER_56_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4530_ _8438_/Q _4533_/C vssd1 vssd1 vccd1 vccd1 _4532_/A sky130_fd_sc_hd__and2_1
X_4461_ _4766_/B vssd1 vssd1 vccd1 vccd1 _4759_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_7180_ _7180_/A _7180_/B _7180_/C vssd1 vssd1 vccd1 vccd1 _7205_/A sky130_fd_sc_hd__or3_4
X_6200_ _6200_/A _6200_/B vssd1 vssd1 vccd1 vccd1 _6201_/B sky130_fd_sc_hd__xnor2_1
X_4392_ _6514_/A vssd1 vssd1 vccd1 vccd1 _5180_/A sky130_fd_sc_hd__clkbuf_1
X_6131_ _6132_/A _6132_/B _6132_/C vssd1 vssd1 vccd1 vccd1 _6131_/X sky130_fd_sc_hd__o21a_1
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6062_ _6063_/A _6063_/B vssd1 vssd1 vccd1 vccd1 _6078_/A sky130_fd_sc_hd__and2b_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5013_ _5099_/A _5093_/B _5093_/C vssd1 vssd1 vccd1 vccd1 _5014_/D sky130_fd_sc_hd__or3_1
XFILLER_78_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6964_ _7032_/A _6964_/B _6964_/C vssd1 vssd1 vccd1 vccd1 _7044_/A sky130_fd_sc_hd__or3_1
X_8703_ _8703_/A _4283_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[20] sky130_fd_sc_hd__ebufn_8
XFILLER_81_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6895_ _6897_/A _6897_/B vssd1 vssd1 vccd1 vccd1 _6895_/Y sky130_fd_sc_hd__nand2_1
X_5915_ _5915_/A _5915_/B vssd1 vssd1 vccd1 vccd1 _5959_/A sky130_fd_sc_hd__xnor2_1
XFILLER_21_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5846_ _5846_/A _6021_/A vssd1 vssd1 vccd1 vccd1 _5846_/Y sky130_fd_sc_hd__nor2_1
X_8565_ input3/X _8565_/D vssd1 vssd1 vccd1 vccd1 _8565_/Q sky130_fd_sc_hd__dfxtp_1
X_5777_ _5825_/A _5838_/A vssd1 vssd1 vccd1 vccd1 _5942_/B sky130_fd_sc_hd__or2_2
X_8496_ input3/X _8496_/D vssd1 vssd1 vccd1 vccd1 _8496_/Q sky130_fd_sc_hd__dfxtp_1
X_4728_ _4766_/C vssd1 vssd1 vccd1 vccd1 _4790_/B sky130_fd_sc_hd__buf_2
XFILLER_5_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7516_ _7505_/A _7505_/B _7507_/X _7508_/A vssd1 vssd1 vccd1 vccd1 _7520_/A sky130_fd_sc_hd__a31o_1
X_4659_ _4659_/A _4659_/B _5179_/B _4659_/D vssd1 vssd1 vccd1 vccd1 _4663_/B sky130_fd_sc_hd__or4_2
X_7447_ _7462_/A vssd1 vssd1 vccd1 vccd1 _8430_/A sky130_fd_sc_hd__buf_2
X_7378_ _7378_/A vssd1 vssd1 vccd1 vccd1 _8561_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6329_ _6382_/B vssd1 vssd1 vccd1 vccd1 _6331_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5700_ _5662_/A _5662_/B _5699_/X vssd1 vssd1 vccd1 vccd1 _5748_/B sky130_fd_sc_hd__o21ai_1
X_6680_ _6680_/A vssd1 vssd1 vccd1 vccd1 _7323_/A sky130_fd_sc_hd__clkbuf_1
X_5631_ _5631_/A _5631_/B _5631_/C vssd1 vssd1 vccd1 vccd1 _5632_/B sky130_fd_sc_hd__nand3_1
X_8350_ _8345_/X _8346_/X _8348_/X _8349_/Y vssd1 vssd1 vccd1 vccd1 _8351_/B sky130_fd_sc_hd__a31oi_2
X_5562_ _5562_/A _5900_/A vssd1 vssd1 vccd1 vccd1 _5578_/A sky130_fd_sc_hd__nand2_1
X_4513_ _6427_/A _8453_/Q vssd1 vssd1 vccd1 vccd1 _4536_/A sky130_fd_sc_hd__nor2_1
X_7301_ _7301_/A _7301_/B vssd1 vssd1 vccd1 vccd1 _7302_/B sky130_fd_sc_hd__xnor2_1
X_8281_ _8281_/A _8281_/B vssd1 vssd1 vccd1 vccd1 _8284_/A sky130_fd_sc_hd__xor2_1
X_7232_ _7232_/A _7232_/B vssd1 vssd1 vccd1 vccd1 _7233_/C sky130_fd_sc_hd__xnor2_1
X_5493_ _5493_/A vssd1 vssd1 vccd1 vccd1 _5499_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4444_ _4670_/A _4706_/B _4470_/A _4464_/C vssd1 vssd1 vccd1 vccd1 _4445_/A sky130_fd_sc_hd__or4_4
X_7163_ _7162_/A _7163_/B vssd1 vssd1 vccd1 vccd1 _7163_/X sky130_fd_sc_hd__and2b_1
X_4375_ _4375_/A vssd1 vssd1 vccd1 vccd1 _4375_/Y sky130_fd_sc_hd__inv_2
X_7094_ _7272_/B _7028_/C _7146_/A vssd1 vssd1 vccd1 vccd1 _7095_/B sky130_fd_sc_hd__a21o_1
X_6114_ _6114_/A _6114_/B vssd1 vssd1 vccd1 vccd1 _6117_/A sky130_fd_sc_hd__xnor2_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6045_ _6098_/A _6045_/B vssd1 vssd1 vccd1 vccd1 _6046_/B sky130_fd_sc_hd__xnor2_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7996_ _7996_/A _8019_/B vssd1 vssd1 vccd1 vccd1 _8013_/A sky130_fd_sc_hd__xnor2_1
X_6947_ _6947_/A _6948_/A _6947_/C vssd1 vssd1 vccd1 vccd1 _7015_/A sky130_fd_sc_hd__or3_2
X_6878_ _6880_/A _6880_/B _6880_/C vssd1 vssd1 vccd1 vccd1 _6878_/X sky130_fd_sc_hd__and3_1
X_5829_ _6025_/B _5829_/B _5829_/C vssd1 vssd1 vccd1 vccd1 _6019_/A sky130_fd_sc_hd__and3b_1
X_8548_ input3/X _8548_/D vssd1 vssd1 vccd1 vccd1 _8548_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8479_ input3/X _8479_/D vssd1 vssd1 vccd1 vccd1 _8479_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7850_ _7888_/B vssd1 vssd1 vccd1 vccd1 _8147_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_63_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6801_ _6802_/B _6802_/C _6980_/B vssd1 vssd1 vccd1 vccd1 _6863_/C sky130_fd_sc_hd__a21o_1
XFILLER_51_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4993_ _4993_/A _4993_/B _4945_/B vssd1 vssd1 vccd1 vccd1 _5169_/B sky130_fd_sc_hd__or3b_2
X_7781_ _7781_/A _7781_/B vssd1 vssd1 vccd1 vccd1 _7786_/A sky130_fd_sc_hd__xnor2_1
X_6732_ _6907_/A _6907_/B _6731_/X vssd1 vssd1 vccd1 vccd1 _6912_/A sky130_fd_sc_hd__o21ai_1
XFILLER_51_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6663_ _6663_/A _6663_/B vssd1 vssd1 vccd1 vccd1 _6663_/Y sky130_fd_sc_hd__nand2_1
X_5614_ _5738_/A _6025_/A vssd1 vssd1 vccd1 vccd1 _5619_/A sky130_fd_sc_hd__nor2_1
X_8402_ _8401_/X _8397_/B _8418_/S vssd1 vssd1 vccd1 vccd1 _8403_/B sky130_fd_sc_hd__mux2_1
X_6594_ _6964_/B vssd1 vssd1 vccd1 vccd1 _7039_/B sky130_fd_sc_hd__clkbuf_2
X_8333_ _8333_/A _8333_/B vssd1 vssd1 vccd1 vccd1 _8337_/A sky130_fd_sc_hd__xnor2_1
X_5545_ _5649_/A _5596_/C vssd1 vssd1 vccd1 vccd1 _5547_/B sky130_fd_sc_hd__xnor2_1
X_8264_ _8264_/A _8264_/B vssd1 vssd1 vccd1 vccd1 _8266_/B sky130_fd_sc_hd__xnor2_1
XFILLER_2_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5476_ _5767_/A _5764_/A vssd1 vssd1 vccd1 vccd1 _5932_/A sky130_fd_sc_hd__or2_1
X_7215_ _7218_/B _7218_/A vssd1 vssd1 vccd1 vccd1 _7215_/X sky130_fd_sc_hd__and2b_1
X_4427_ _8467_/Q vssd1 vssd1 vccd1 vccd1 _7494_/B sky130_fd_sc_hd__clkbuf_4
X_8195_ _8196_/A _8196_/B vssd1 vssd1 vccd1 vccd1 _8207_/B sky130_fd_sc_hd__xnor2_1
X_7146_ _7146_/A _7146_/B _7146_/C vssd1 vssd1 vccd1 vccd1 _7345_/A sky130_fd_sc_hd__and3_1
X_4358_ _4358_/A vssd1 vssd1 vccd1 vccd1 _4363_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_48_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4289_ _4289_/A vssd1 vssd1 vccd1 vccd1 _4289_/Y sky130_fd_sc_hd__inv_2
X_7077_ _7077_/A _7077_/B vssd1 vssd1 vccd1 vccd1 _7077_/Y sky130_fd_sc_hd__nor2_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8671__87 vssd1 vssd1 vccd1 vccd1 _8671__87/HI _8780_/A sky130_fd_sc_hd__conb_1
XFILLER_27_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6028_ _6135_/A _6135_/B vssd1 vssd1 vccd1 vccd1 _6030_/A sky130_fd_sc_hd__xnor2_2
XFILLER_27_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7979_ _8024_/A vssd1 vssd1 vccd1 vccd1 _8120_/A sky130_fd_sc_hd__inv_2
XFILLER_42_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_80 _8789_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5330_ _5332_/A _5333_/A _5374_/A vssd1 vssd1 vccd1 vccd1 _5331_/A sky130_fd_sc_hd__mux2_1
X_5261_ _5263_/B _5261_/B _5294_/A vssd1 vssd1 vccd1 vccd1 _5262_/A sky130_fd_sc_hd__and3b_1
XFILLER_5_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7000_ _7002_/A vssd1 vssd1 vccd1 vccd1 _7248_/A sky130_fd_sc_hd__clkbuf_2
X_5192_ _8475_/Q _5192_/B vssd1 vssd1 vccd1 vccd1 _5192_/X sky130_fd_sc_hd__or2_1
XFILLER_68_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7902_ _7902_/A _7902_/B vssd1 vssd1 vccd1 vccd1 _7903_/B sky130_fd_sc_hd__xnor2_4
XFILLER_91_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7833_ _7834_/A _7834_/B vssd1 vssd1 vccd1 vccd1 _8012_/A sky130_fd_sc_hd__nand2_1
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7764_ _7695_/B _7763_/Y _7652_/B _7658_/B vssd1 vssd1 vccd1 vccd1 _7802_/A sky130_fd_sc_hd__a22o_1
X_4976_ _4976_/A _5088_/B _5022_/B vssd1 vssd1 vccd1 vccd1 _5009_/C sky130_fd_sc_hd__or3_1
X_6715_ _6941_/A _6715_/B vssd1 vssd1 vccd1 vccd1 _6987_/B sky130_fd_sc_hd__xnor2_4
X_7695_ _7804_/A _7695_/B vssd1 vssd1 vccd1 vccd1 _7697_/A sky130_fd_sc_hd__nand2_1
X_6646_ _6896_/B _6896_/C _6896_/A vssd1 vssd1 vccd1 vccd1 _6663_/A sky130_fd_sc_hd__a21bo_1
X_6577_ _6683_/A _6683_/B vssd1 vssd1 vccd1 vccd1 _7069_/B sky130_fd_sc_hd__or2_2
X_8316_ _8269_/A _8269_/B _8267_/A vssd1 vssd1 vccd1 vccd1 _8333_/A sky130_fd_sc_hd__o21a_1
X_5528_ _5703_/A _5528_/B vssd1 vssd1 vccd1 vccd1 _5530_/A sky130_fd_sc_hd__nand2_1
XFILLER_3_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8247_ _8247_/A _8247_/B vssd1 vssd1 vccd1 vccd1 _8255_/A sky130_fd_sc_hd__nor2_1
X_5459_ _5459_/A _5459_/B vssd1 vssd1 vccd1 vccd1 _5492_/B sky130_fd_sc_hd__xnor2_4
X_8178_ _8198_/A _8198_/B vssd1 vssd1 vccd1 vccd1 _8194_/A sky130_fd_sc_hd__xor2_1
X_7129_ _7129_/A _7129_/B vssd1 vssd1 vccd1 vccd1 _7129_/X sky130_fd_sc_hd__or2_1
XFILLER_59_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4830_ _5151_/C _5147_/B _5018_/A vssd1 vssd1 vccd1 vccd1 _4830_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_33_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4761_ _8465_/Q _4761_/B _4766_/C vssd1 vssd1 vccd1 vccd1 _4791_/A sky130_fd_sc_hd__or3_4
X_6500_ _6500_/A _6500_/B vssd1 vssd1 vccd1 vccd1 _6534_/A sky130_fd_sc_hd__xnor2_2
X_4692_ _4692_/A vssd1 vssd1 vccd1 vccd1 _8469_/D sky130_fd_sc_hd__clkbuf_1
X_7480_ _7477_/A _7477_/C _7477_/B vssd1 vssd1 vccd1 vccd1 _7484_/A sky130_fd_sc_hd__a21bo_1
X_6431_ _6431_/A vssd1 vssd1 vccd1 vccd1 _8550_/D sky130_fd_sc_hd__clkbuf_1
X_6362_ _8538_/Q _6362_/B _6362_/C vssd1 vssd1 vccd1 vccd1 _6366_/B sky130_fd_sc_hd__and3_1
X_8101_ _8041_/A _8229_/A _8101_/C vssd1 vssd1 vccd1 vccd1 _8229_/B sky130_fd_sc_hd__nand3b_1
X_5313_ _8513_/Q vssd1 vssd1 vccd1 vccd1 _5366_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6293_ _6293_/A _6293_/B vssd1 vssd1 vccd1 vccd1 _6297_/B sky130_fd_sc_hd__nor2_1
XFILLER_88_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5244_ _6396_/B _5246_/C _5230_/B vssd1 vssd1 vccd1 vccd1 _5244_/Y sky130_fd_sc_hd__o21ai_1
X_8032_ _7827_/X _8005_/B _8003_/Y vssd1 vssd1 vccd1 vccd1 _8034_/B sky130_fd_sc_hd__a21oi_2
X_5175_ _5158_/X _5174_/X _5175_/S vssd1 vssd1 vccd1 vccd1 _5175_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8641__57 vssd1 vssd1 vccd1 vccd1 _8641__57/HI _8750_/A sky130_fd_sc_hd__conb_1
XFILLER_36_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7816_ _7817_/A _7817_/B vssd1 vssd1 vccd1 vccd1 _7933_/B sky130_fd_sc_hd__or2_1
XFILLER_36_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4959_ _4955_/X _4957_/X _4991_/A _5117_/A vssd1 vssd1 vccd1 vccd1 _4959_/X sky130_fd_sc_hd__a211o_1
XFILLER_61_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7747_ _7747_/A _7945_/A vssd1 vssd1 vccd1 vccd1 _7748_/B sky130_fd_sc_hd__nand2_1
XFILLER_20_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7678_ _7678_/A _7678_/B vssd1 vssd1 vccd1 vccd1 _7690_/A sky130_fd_sc_hd__or2_1
X_6629_ _6969_/B _6969_/C vssd1 vssd1 vccd1 vccd1 _7043_/B sky130_fd_sc_hd__nand2_2
XFILLER_10_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6980_ _6980_/A _6980_/B vssd1 vssd1 vccd1 vccd1 _6981_/S sky130_fd_sc_hd__nand2_1
XFILLER_26_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5931_ _5826_/A _5930_/Y _6243_/B vssd1 vssd1 vccd1 vccd1 _6200_/A sky130_fd_sc_hd__o21a_1
X_5862_ _5859_/B _5860_/Y _5861_/X vssd1 vssd1 vccd1 vccd1 _5863_/B sky130_fd_sc_hd__a21boi_1
X_4813_ _4953_/A _4944_/A _4786_/B vssd1 vssd1 vccd1 vccd1 _4869_/B sky130_fd_sc_hd__a21oi_1
X_5793_ _5793_/A _6108_/A vssd1 vssd1 vccd1 vccd1 _6226_/A sky130_fd_sc_hd__xor2_4
XFILLER_21_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7601_ _7612_/A _7616_/B vssd1 vssd1 vccd1 vccd1 _7604_/A sky130_fd_sc_hd__nand2_2
X_8581_ input3/X _8581_/D vssd1 vssd1 vccd1 vccd1 _8581_/Q sky130_fd_sc_hd__dfxtp_1
X_4744_ _4805_/A _4818_/B vssd1 vssd1 vccd1 vccd1 _5160_/C sky130_fd_sc_hd__nor2_2
X_7532_ _7679_/A _7532_/B vssd1 vssd1 vccd1 vccd1 _7682_/B sky130_fd_sc_hd__xnor2_1
X_4675_ _4790_/A _4675_/B vssd1 vssd1 vccd1 vccd1 _4676_/A sky130_fd_sc_hd__or2_1
X_7463_ _7461_/Y _7501_/A _8418_/S vssd1 vssd1 vccd1 vccd1 _7464_/B sky130_fd_sc_hd__mux2_1
X_7394_ _6562_/B _5241_/X _6432_/A _7393_/X vssd1 vssd1 vccd1 vccd1 _8564_/D sky130_fd_sc_hd__a22o_1
X_6414_ _8551_/Q vssd1 vssd1 vccd1 vccd1 _6433_/A sky130_fd_sc_hd__clkbuf_2
X_6345_ _6351_/C _6345_/B _6382_/B vssd1 vssd1 vccd1 vccd1 _6346_/A sky130_fd_sc_hd__and3b_1
X_6276_ _6276_/A _6276_/B vssd1 vssd1 vccd1 vccd1 _6278_/A sky130_fd_sc_hd__nor2_1
XFILLER_88_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5227_ _8505_/Q _8504_/Q _5226_/X _8506_/Q vssd1 vssd1 vccd1 vccd1 _6465_/A sky130_fd_sc_hd__a31oi_4
X_8015_ _8015_/A _8015_/B _7872_/B vssd1 vssd1 vccd1 vccd1 _8188_/A sky130_fd_sc_hd__or3b_1
XFILLER_88_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5158_ _5174_/S _4943_/B _5152_/X _5157_/X _4623_/X vssd1 vssd1 vccd1 vccd1 _5158_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_29_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5089_ _5089_/A _5089_/B _5089_/C _5089_/D vssd1 vssd1 vccd1 vccd1 _5089_/X sky130_fd_sc_hd__or4_1
XFILLER_84_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8779_ _8779_/A _4373_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[26] sky130_fd_sc_hd__ebufn_8
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4460_ _8464_/Q vssd1 vssd1 vccd1 vccd1 _4766_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_4391_ _8462_/Q vssd1 vssd1 vccd1 vccd1 _6514_/A sky130_fd_sc_hd__clkbuf_4
X_6130_ _6193_/A _6130_/B vssd1 vssd1 vccd1 vccd1 _6132_/C sky130_fd_sc_hd__nand2_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6061_ _6061_/A _6061_/B vssd1 vssd1 vccd1 vccd1 _6063_/B sky130_fd_sc_hd__xor2_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5012_ _5012_/A _5055_/B _5012_/C _5028_/D vssd1 vssd1 vccd1 vccd1 _5012_/X sky130_fd_sc_hd__or4_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8611__27 vssd1 vssd1 vccd1 vccd1 _8611__27/HI _8706_/A sky130_fd_sc_hd__conb_1
XFILLER_38_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6963_ _7093_/A _6963_/B vssd1 vssd1 vccd1 vccd1 _7272_/A sky130_fd_sc_hd__xnor2_1
XFILLER_81_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8702_ _8702_/A _4282_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[19] sky130_fd_sc_hd__ebufn_8
X_6894_ _7297_/A _6894_/B vssd1 vssd1 vccd1 vccd1 _6897_/B sky130_fd_sc_hd__xor2_2
XFILLER_53_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5914_ _5914_/A _5914_/B vssd1 vssd1 vccd1 vccd1 _5915_/B sky130_fd_sc_hd__nand2_1
XFILLER_34_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5845_ _5925_/A _5925_/B vssd1 vssd1 vccd1 vccd1 _5853_/A sky130_fd_sc_hd__xor2_2
XFILLER_34_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8564_ input3/X _8564_/D vssd1 vssd1 vccd1 vccd1 _8564_/Q sky130_fd_sc_hd__dfxtp_1
X_5776_ _5776_/A _5776_/B vssd1 vssd1 vccd1 vccd1 _5823_/A sky130_fd_sc_hd__and2_2
X_8495_ input3/X _8495_/D vssd1 vssd1 vccd1 vccd1 _8495_/Q sky130_fd_sc_hd__dfxtp_1
X_4727_ _7494_/B _8466_/Q vssd1 vssd1 vccd1 vccd1 _4766_/C sky130_fd_sc_hd__or2_1
X_7515_ _7804_/A _8367_/B vssd1 vssd1 vccd1 vccd1 _7530_/A sky130_fd_sc_hd__nand2_1
X_4658_ _4658_/A vssd1 vssd1 vccd1 vccd1 _8463_/D sky130_fd_sc_hd__clkbuf_1
X_7446_ _8570_/Q vssd1 vssd1 vccd1 vccd1 _7494_/A sky130_fd_sc_hd__inv_2
XFILLER_89_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7377_ _5294_/A _6428_/A _7377_/S vssd1 vssd1 vccd1 vccd1 _7378_/A sky130_fd_sc_hd__mux2_1
X_4589_ _4762_/C vssd1 vssd1 vccd1 vccd1 _4675_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6328_ _6328_/A _6328_/B vssd1 vssd1 vccd1 vccd1 _6382_/B sky130_fd_sc_hd__and2_2
XFILLER_88_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6259_ _6259_/A _6259_/B vssd1 vssd1 vccd1 vccd1 _6259_/Y sky130_fd_sc_hd__nand2_1
XFILLER_88_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8677__93 vssd1 vssd1 vccd1 vccd1 _8677__93/HI _8786_/A sky130_fd_sc_hd__conb_1
XFILLER_95_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5630_ _5631_/A _5631_/B _5631_/C vssd1 vssd1 vccd1 vccd1 _5719_/A sky130_fd_sc_hd__a21o_1
X_5561_ _5561_/A _5561_/B vssd1 vssd1 vccd1 vccd1 _5574_/A sky130_fd_sc_hd__or2_1
X_4512_ input2/X vssd1 vssd1 vccd1 vccd1 _6427_/A sky130_fd_sc_hd__inv_2
X_7300_ _7300_/A _7300_/B vssd1 vssd1 vccd1 vccd1 _7301_/B sky130_fd_sc_hd__xnor2_1
X_8280_ _8334_/A _8334_/B vssd1 vssd1 vccd1 vccd1 _8281_/B sky130_fd_sc_hd__xnor2_1
X_5492_ _5615_/A _5492_/B vssd1 vssd1 vccd1 vccd1 _5502_/A sky130_fd_sc_hd__nor2_1
X_7231_ _7228_/B _7228_/C _7228_/A vssd1 vssd1 vccd1 vccd1 _7241_/B sky130_fd_sc_hd__o21ai_1
X_4443_ _7766_/B _4706_/A vssd1 vssd1 vccd1 vccd1 _4464_/C sky130_fd_sc_hd__nand2_1
X_7162_ _7162_/A _7163_/B vssd1 vssd1 vccd1 vccd1 _7194_/B sky130_fd_sc_hd__xnor2_1
X_4374_ _4375_/A vssd1 vssd1 vccd1 vccd1 _4374_/Y sky130_fd_sc_hd__inv_2
X_7093_ _7093_/A _7098_/B _7093_/C vssd1 vssd1 vccd1 vccd1 _7264_/A sky130_fd_sc_hd__nor3_1
X_6113_ _6211_/A _6211_/B vssd1 vssd1 vccd1 vccd1 _6114_/B sky130_fd_sc_hd__xor2_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6044_ _6044_/A _6044_/B vssd1 vssd1 vccd1 vccd1 _6045_/B sky130_fd_sc_hd__xnor2_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8592__8 vssd1 vssd1 vccd1 vccd1 _8592__8/HI _8687_/A sky130_fd_sc_hd__conb_1
XFILLER_93_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7995_ _7995_/A _7995_/B vssd1 vssd1 vccd1 vccd1 _8019_/B sky130_fd_sc_hd__xor2_1
X_6946_ _6945_/A _6945_/C _6945_/B vssd1 vssd1 vccd1 vccd1 _6947_/C sky130_fd_sc_hd__a21oi_1
X_6877_ _6874_/B _6874_/C _6812_/A vssd1 vssd1 vccd1 vccd1 _6880_/C sky130_fd_sc_hd__a21o_1
XFILLER_22_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5828_ _5828_/A _6137_/A vssd1 vssd1 vccd1 vccd1 _5829_/B sky130_fd_sc_hd__nand2_1
X_8547_ input3/X _8547_/D vssd1 vssd1 vccd1 vccd1 _8547_/Q sky130_fd_sc_hd__dfxtp_1
X_5759_ _5757_/X _5735_/B _5758_/Y vssd1 vssd1 vccd1 vccd1 _5821_/A sky130_fd_sc_hd__a21bo_2
X_8478_ input3/X _8478_/D vssd1 vssd1 vccd1 vccd1 _8478_/Q sky130_fd_sc_hd__dfxtp_1
X_7429_ _7416_/X _7417_/A _8423_/B vssd1 vssd1 vccd1 vccd1 _7429_/X sky130_fd_sc_hd__a21bo_1
XFILLER_89_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6800_ _6980_/A _7291_/B _7291_/A vssd1 vssd1 vccd1 vccd1 _6863_/B sky130_fd_sc_hd__a21o_1
X_4992_ _5039_/B _5053_/B _5018_/C _4992_/D vssd1 vssd1 vccd1 vccd1 _4992_/X sky130_fd_sc_hd__or4_1
XFILLER_63_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7780_ _7804_/C _7780_/B vssd1 vssd1 vccd1 vccd1 _7781_/B sky130_fd_sc_hd__xnor2_1
X_6731_ _6731_/A _6731_/B vssd1 vssd1 vccd1 vccd1 _6731_/X sky130_fd_sc_hd__or2_1
XFILLER_23_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6662_ _6663_/A _6663_/B vssd1 vssd1 vccd1 vccd1 _6902_/B sky130_fd_sc_hd__xnor2_1
X_5613_ _5722_/B _5612_/C _5612_/A vssd1 vssd1 vccd1 vccd1 _5620_/B sky130_fd_sc_hd__a21oi_1
X_8401_ _8401_/A _8401_/B vssd1 vssd1 vccd1 vccd1 _8401_/X sky130_fd_sc_hd__xor2_1
X_6593_ _6614_/A vssd1 vssd1 vccd1 vccd1 _6964_/B sky130_fd_sc_hd__clkbuf_2
X_8332_ _8332_/A _8332_/B vssd1 vssd1 vccd1 vccd1 _8333_/B sky130_fd_sc_hd__xnor2_1
X_5544_ _5664_/A _5544_/B vssd1 vssd1 vccd1 vccd1 _5596_/C sky130_fd_sc_hd__xnor2_1
X_8263_ _8263_/A _8321_/B vssd1 vssd1 vccd1 vccd1 _8264_/B sky130_fd_sc_hd__xnor2_1
X_5475_ _5492_/B vssd1 vssd1 vccd1 vccd1 _5764_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7214_ _7152_/A _7148_/B _7005_/X vssd1 vssd1 vccd1 vccd1 _7218_/A sky130_fd_sc_hd__o21ai_1
X_4426_ _4698_/A _4466_/B _4715_/A vssd1 vssd1 vccd1 vccd1 _4464_/B sky130_fd_sc_hd__nand3_1
X_8194_ _8194_/A _8194_/B vssd1 vssd1 vccd1 vccd1 _8196_/B sky130_fd_sc_hd__xnor2_1
X_7145_ _7143_/X _7142_/Y _7141_/X _7137_/X vssd1 vssd1 vccd1 vccd1 _7146_/C sky130_fd_sc_hd__a211o_1
XFILLER_86_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4357_ _4357_/A vssd1 vssd1 vccd1 vccd1 _4357_/Y sky130_fd_sc_hd__inv_2
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4288_ _4289_/A vssd1 vssd1 vccd1 vccd1 _4288_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7076_ _7131_/A _7131_/B vssd1 vssd1 vccd1 vccd1 _7081_/A sky130_fd_sc_hd__nand2_1
XFILLER_86_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6027_ _6137_/C _6027_/B vssd1 vssd1 vccd1 vccd1 _6135_/B sky130_fd_sc_hd__xnor2_1
XFILLER_27_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7978_ _7978_/A _7978_/B vssd1 vssd1 vccd1 vccd1 _8024_/A sky130_fd_sc_hd__or2_1
X_6929_ _6929_/A _6929_/B vssd1 vssd1 vccd1 vccd1 _6930_/B sky130_fd_sc_hd__or2_1
XFILLER_22_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8647__63 vssd1 vssd1 vccd1 vccd1 _8647__63/HI _8756_/A sky130_fd_sc_hd__conb_1
XFILLER_49_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_70 _8783_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_81 _8789_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5260_ _5260_/A vssd1 vssd1 vccd1 vccd1 _5294_/A sky130_fd_sc_hd__buf_2
XFILLER_5_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5191_ _8516_/Q _5188_/X _5189_/X _6426_/A vssd1 vssd1 vccd1 vccd1 _8474_/D sky130_fd_sc_hd__o211a_1
XFILLER_55_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7901_ _7944_/A _7901_/B vssd1 vssd1 vccd1 vccd1 _7902_/B sky130_fd_sc_hd__xor2_4
X_7832_ _8037_/A _7832_/B vssd1 vssd1 vccd1 vccd1 _7834_/B sky130_fd_sc_hd__nor2_1
X_4975_ _5171_/B _4975_/B _4975_/C vssd1 vssd1 vccd1 vccd1 _5022_/B sky130_fd_sc_hd__or3_2
XFILLER_51_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7763_ _7824_/A _8097_/A vssd1 vssd1 vccd1 vccd1 _7763_/Y sky130_fd_sc_hd__nor2_1
X_6714_ _6714_/A _6714_/B _6714_/C vssd1 vssd1 vccd1 vccd1 _6715_/B sky130_fd_sc_hd__or3_2
X_7694_ _7694_/A _7694_/B vssd1 vssd1 vccd1 vccd1 _8371_/A sky130_fd_sc_hd__xnor2_2
X_6645_ _6645_/A _6733_/B _6645_/C vssd1 vssd1 vccd1 vccd1 _6896_/A sky130_fd_sc_hd__nand3_1
XFILLER_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6576_ _6575_/B _6575_/C _6575_/A vssd1 vssd1 vccd1 vccd1 _6683_/B sky130_fd_sc_hd__a21oi_1
X_8315_ _8315_/A _8315_/B vssd1 vssd1 vccd1 vccd1 _8343_/A sky130_fd_sc_hd__xnor2_1
X_5527_ _8515_/Q _7644_/B vssd1 vssd1 vccd1 vccd1 _5528_/B sky130_fd_sc_hd__nand2_1
X_8246_ _8167_/A _8166_/B _8166_/A vssd1 vssd1 vccd1 vccd1 _8286_/A sky130_fd_sc_hd__o21ba_1
XFILLER_59_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5458_ _5828_/A vssd1 vssd1 vccd1 vccd1 _5846_/A sky130_fd_sc_hd__clkbuf_2
X_4409_ _8466_/Q vssd1 vssd1 vccd1 vccd1 _4718_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5389_ _5563_/A _5563_/B vssd1 vssd1 vccd1 vccd1 _5800_/A sky130_fd_sc_hd__xnor2_4
X_8177_ _7834_/A _8176_/Y _7804_/C _7780_/B vssd1 vssd1 vccd1 vccd1 _8198_/B sky130_fd_sc_hd__a2bb2o_1
X_7128_ _7151_/A _7151_/B vssd1 vssd1 vccd1 vccd1 _7133_/A sky130_fd_sc_hd__nor2_1
XFILLER_59_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7059_ _7077_/A _7077_/B vssd1 vssd1 vccd1 vccd1 _7060_/B sky130_fd_sc_hd__xor2_1
XFILLER_46_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4760_ _4779_/A _4792_/A vssd1 vssd1 vccd1 vccd1 _4760_/Y sky130_fd_sc_hd__nor2_1
XFILLER_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4691_ _4698_/C _7412_/A _4691_/C vssd1 vssd1 vccd1 vccd1 _4692_/A sky130_fd_sc_hd__and3b_1
X_6430_ _5294_/A _6432_/A _6435_/A vssd1 vssd1 vccd1 vccd1 _6431_/A sky130_fd_sc_hd__mux2_1
X_6361_ _6362_/B _6362_/C _6360_/Y vssd1 vssd1 vccd1 vccd1 _8537_/D sky130_fd_sc_hd__a21oi_1
X_8100_ _8101_/C _8229_/A _7695_/B vssd1 vssd1 vccd1 vccd1 _8102_/B sky130_fd_sc_hd__a21o_1
X_5312_ _8514_/Q vssd1 vssd1 vccd1 vccd1 _5360_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6292_ _6293_/A _6293_/B vssd1 vssd1 vccd1 vccd1 _6294_/A sky130_fd_sc_hd__and2_1
X_5243_ _5246_/C _5243_/B vssd1 vssd1 vccd1 vccd1 _8489_/D sky130_fd_sc_hd__nor2_1
X_8031_ _8092_/A _8031_/B vssd1 vssd1 vccd1 vccd1 _8034_/A sky130_fd_sc_hd__xnor2_2
X_5174_ _5166_/X _5173_/X _5174_/S vssd1 vssd1 vccd1 vccd1 _5174_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7815_ _7830_/B _7815_/B vssd1 vssd1 vccd1 vccd1 _7817_/B sky130_fd_sc_hd__xnor2_1
XFILLER_51_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4958_ _4970_/A vssd1 vssd1 vccd1 vccd1 _5117_/A sky130_fd_sc_hd__clkbuf_2
X_7746_ _7746_/A vssd1 vssd1 vccd1 vccd1 _7945_/A sky130_fd_sc_hd__clkbuf_2
X_4889_ _5019_/B _4975_/B vssd1 vssd1 vccd1 vccd1 _4890_/A sky130_fd_sc_hd__nor2_1
X_7677_ _7677_/A _7677_/B vssd1 vssd1 vccd1 vccd1 _7678_/B sky130_fd_sc_hd__and2_1
X_6628_ _6627_/B _6627_/C _6627_/A vssd1 vssd1 vccd1 vccd1 _6969_/C sky130_fd_sc_hd__a21o_1
XFILLER_20_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6559_ _6939_/A _6941_/A vssd1 vssd1 vccd1 vccd1 _6560_/B sky130_fd_sc_hd__nor2_1
XFILLER_79_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8229_ _8229_/A _8229_/B vssd1 vssd1 vccd1 vccd1 _8235_/A sky130_fd_sc_hd__nand2_1
XFILLER_86_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8617__33 vssd1 vssd1 vccd1 vccd1 _8617__33/HI _8712_/A sky130_fd_sc_hd__conb_1
XFILLER_59_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5930_ _5930_/A _5930_/B vssd1 vssd1 vccd1 vccd1 _5930_/Y sky130_fd_sc_hd__nor2_1
XFILLER_34_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5861_ _5861_/A _5984_/A _5861_/C vssd1 vssd1 vccd1 vccd1 _5861_/X sky130_fd_sc_hd__or3_1
X_7600_ _8586_/Q _8462_/Q vssd1 vssd1 vccd1 vccd1 _7616_/B sky130_fd_sc_hd__or2b_1
X_4812_ _4812_/A vssd1 vssd1 vccd1 vccd1 _4944_/A sky130_fd_sc_hd__inv_2
X_8580_ input3/X _8580_/D vssd1 vssd1 vccd1 vccd1 _8580_/Q sky130_fd_sc_hd__dfxtp_1
X_5792_ _5792_/A vssd1 vssd1 vccd1 vccd1 _6108_/A sky130_fd_sc_hd__buf_2
XFILLER_21_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4743_ _4796_/B vssd1 vssd1 vccd1 vccd1 _4818_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_21_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7531_ _7824_/A _7530_/A _7983_/A _7530_/Y vssd1 vssd1 vccd1 vccd1 _7532_/B sky130_fd_sc_hd__o31a_1
X_7462_ _7462_/A vssd1 vssd1 vccd1 vccd1 _8418_/S sky130_fd_sc_hd__buf_2
X_6413_ _8555_/Q vssd1 vssd1 vccd1 vccd1 _6541_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4674_ _4689_/A vssd1 vssd1 vccd1 vccd1 _8403_/A sky130_fd_sc_hd__buf_2
X_7393_ _7393_/A _7393_/B vssd1 vssd1 vccd1 vccd1 _7393_/X sky130_fd_sc_hd__xor2_1
X_6344_ _8530_/Q _6319_/D _6338_/B _8532_/Q vssd1 vssd1 vccd1 vccd1 _6345_/B sky130_fd_sc_hd__a31o_1
XFILLER_88_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6275_ _6274_/B _6281_/B vssd1 vssd1 vccd1 vccd1 _6276_/B sky130_fd_sc_hd__and2b_1
X_5226_ _8503_/Q _8502_/Q _5226_/C vssd1 vssd1 vccd1 vccd1 _5226_/X sky130_fd_sc_hd__or3_1
X_8014_ _8016_/A _8016_/B vssd1 vssd1 vccd1 vccd1 _8190_/A sky130_fd_sc_hd__and2_1
X_5157_ _4947_/C _5154_/X _5147_/X _5156_/X vssd1 vssd1 vccd1 vccd1 _5157_/X sky130_fd_sc_hd__o31a_1
XFILLER_56_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5088_ _5088_/A _5088_/B _5088_/C vssd1 vssd1 vccd1 vccd1 _5089_/D sky130_fd_sc_hd__or3_1
XFILLER_84_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8778_ _8778_/A _4372_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[25] sky130_fd_sc_hd__ebufn_8
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7729_ _7841_/B _7728_/C _7728_/A vssd1 vssd1 vccd1 vccd1 _7736_/B sky130_fd_sc_hd__a21oi_1
XFILLER_21_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4390_ _4390_/A vssd1 vssd1 vccd1 vccd1 _4390_/Y sky130_fd_sc_hd__inv_2
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6060_ _6071_/A _6071_/B _6059_/X vssd1 vssd1 vccd1 vccd1 _6063_/A sky130_fd_sc_hd__a21oi_1
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5011_ _5011_/A _5093_/C vssd1 vssd1 vccd1 vccd1 _5092_/D sky130_fd_sc_hd__or2_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6962_ _6962_/A _6962_/B vssd1 vssd1 vccd1 vccd1 _6963_/B sky130_fd_sc_hd__xnor2_1
XFILLER_81_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8701_ _8701_/A _4281_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[18] sky130_fd_sc_hd__ebufn_8
X_6893_ _6893_/A _6913_/B vssd1 vssd1 vccd1 vccd1 _6897_/A sky130_fd_sc_hd__and2_1
XFILLER_53_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5913_ _5965_/A _5965_/B vssd1 vssd1 vccd1 vccd1 _5915_/A sky130_fd_sc_hd__xor2_1
XFILLER_61_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5844_ _5844_/A _5844_/B vssd1 vssd1 vccd1 vccd1 _5925_/B sky130_fd_sc_hd__xnor2_1
XFILLER_22_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8563_ input3/X _8563_/D vssd1 vssd1 vccd1 vccd1 _8563_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5775_ _5739_/A _5767_/X _5740_/B _5826_/A vssd1 vssd1 vccd1 vccd1 _5781_/A sky130_fd_sc_hd__a2bb2o_2
X_7514_ _7768_/A vssd1 vssd1 vccd1 vccd1 _8367_/B sky130_fd_sc_hd__clkbuf_2
X_4726_ _4773_/A _4800_/A vssd1 vssd1 vccd1 vccd1 _5040_/B sky130_fd_sc_hd__nor2_1
X_8494_ input3/X _8494_/D vssd1 vssd1 vccd1 vccd1 _8494_/Q sky130_fd_sc_hd__dfxtp_1
X_4657_ _4657_/A _4657_/B _4657_/C vssd1 vssd1 vccd1 vccd1 _4658_/A sky130_fd_sc_hd__and3_1
X_7445_ _7481_/B _7417_/Y _7442_/Y _7444_/X _6462_/X vssd1 vssd1 vccd1 vccd1 _8569_/D
+ sky130_fd_sc_hd__a221o_1
X_7376_ _8561_/Q vssd1 vssd1 vccd1 vccd1 _7377_/S sky130_fd_sc_hd__inv_2
X_4588_ _4725_/A _4718_/A vssd1 vssd1 vccd1 vccd1 _4762_/C sky130_fd_sc_hd__nand2_1
X_6327_ _6327_/A vssd1 vssd1 vccd1 vccd1 _8527_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6258_ _6259_/A _6259_/B vssd1 vssd1 vccd1 vccd1 _6263_/S sky130_fd_sc_hd__or2_1
X_5209_ _8580_/Q _5202_/X _5208_/X _5200_/X vssd1 vssd1 vccd1 vccd1 _8481_/D sky130_fd_sc_hd__o211a_1
X_6189_ _5839_/A _5618_/A _6188_/Y vssd1 vssd1 vccd1 vccd1 _6189_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_72_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5560_ _5560_/A _5560_/B vssd1 vssd1 vccd1 vccd1 _5561_/B sky130_fd_sc_hd__and2_1
XFILLER_31_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5491_ _5518_/C _5604_/B vssd1 vssd1 vccd1 vccd1 _5504_/A sky130_fd_sc_hd__xnor2_1
X_4511_ _8433_/Q _4511_/B vssd1 vssd1 vccd1 vccd1 _8433_/D sky130_fd_sc_hd__nor2_1
X_7230_ _7256_/A _7256_/B vssd1 vssd1 vccd1 vccd1 _7354_/A sky130_fd_sc_hd__xor2_1
X_4442_ _8472_/Q vssd1 vssd1 vccd1 vccd1 _4706_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7161_ _7161_/A _7161_/B vssd1 vssd1 vccd1 vccd1 _7163_/B sky130_fd_sc_hd__xor2_1
X_4373_ _4375_/A vssd1 vssd1 vccd1 vccd1 _4373_/Y sky130_fd_sc_hd__inv_2
X_7092_ _7090_/X _7089_/Y _7088_/Y _7143_/A vssd1 vssd1 vccd1 vccd1 _7093_/C sky130_fd_sc_hd__a211oi_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6112_ _6112_/A _6112_/B vssd1 vssd1 vccd1 vccd1 _6211_/B sky130_fd_sc_hd__xor2_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6043_ _6043_/A _6043_/B vssd1 vssd1 vccd1 vccd1 _6044_/B sky130_fd_sc_hd__nor2_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7994_ _7994_/A _7994_/B vssd1 vssd1 vccd1 vccd1 _7995_/B sky130_fd_sc_hd__and2_1
X_6945_ _6945_/A _6945_/B _6945_/C vssd1 vssd1 vccd1 vccd1 _6948_/A sky130_fd_sc_hd__and3_1
XFILLER_54_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6876_ _7297_/A _6894_/B vssd1 vssd1 vccd1 vccd1 _6880_/B sky130_fd_sc_hd__nor2_1
XFILLER_10_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5827_ _5940_/A _5827_/B vssd1 vssd1 vccd1 vccd1 _5833_/A sky130_fd_sc_hd__xnor2_2
X_8546_ input3/X _8546_/D vssd1 vssd1 vccd1 vccd1 _8546_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5758_ _5758_/A _5758_/B vssd1 vssd1 vccd1 vccd1 _5758_/Y sky130_fd_sc_hd__nand2_1
X_8477_ input3/X _8477_/D vssd1 vssd1 vccd1 vccd1 _8477_/Q sky130_fd_sc_hd__dfxtp_1
X_4709_ _8410_/A _4709_/B vssd1 vssd1 vccd1 vccd1 _8473_/D sky130_fd_sc_hd__nor2_1
X_5689_ _5689_/A _6118_/A vssd1 vssd1 vccd1 vccd1 _5711_/B sky130_fd_sc_hd__xnor2_2
X_7428_ _7416_/X _7417_/Y _7420_/X _7427_/X vssd1 vssd1 vccd1 vccd1 _7428_/X sky130_fd_sc_hd__o31a_1
X_7359_ _7359_/A _7359_/B vssd1 vssd1 vccd1 vccd1 _7365_/B sky130_fd_sc_hd__and2_1
XFILLER_94_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4991_ _4991_/A _5055_/A _5160_/C _5074_/B vssd1 vssd1 vccd1 vccd1 _4992_/D sky130_fd_sc_hd__or4_1
X_6730_ _6947_/A _6951_/B _6729_/Y vssd1 vssd1 vccd1 vccd1 _6907_/B sky130_fd_sc_hd__o21ba_1
XFILLER_90_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6661_ _6886_/A _6661_/B vssd1 vssd1 vccd1 vccd1 _6663_/B sky130_fd_sc_hd__and2_1
X_6592_ _6592_/A _6592_/B vssd1 vssd1 vccd1 vccd1 _6614_/A sky130_fd_sc_hd__xnor2_1
XFILLER_31_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5612_ _5612_/A _5722_/B _5612_/C vssd1 vssd1 vccd1 vccd1 _5620_/A sky130_fd_sc_hd__and3_1
X_8400_ _8387_/Y _8393_/B _8392_/A vssd1 vssd1 vccd1 vccd1 _8401_/B sky130_fd_sc_hd__o21ai_2
X_8331_ _8331_/A _8331_/B vssd1 vssd1 vccd1 vccd1 _8332_/B sky130_fd_sc_hd__xnor2_1
X_5543_ _5543_/A _5543_/B vssd1 vssd1 vccd1 vccd1 _5544_/B sky130_fd_sc_hd__xor2_1
X_8262_ _7635_/C _7952_/A _8326_/B vssd1 vssd1 vccd1 vccd1 _8321_/B sky130_fd_sc_hd__a21oi_1
X_5474_ _5724_/A vssd1 vssd1 vccd1 vccd1 _6188_/B sky130_fd_sc_hd__buf_2
X_7213_ _7226_/A _7213_/B vssd1 vssd1 vccd1 vccd1 _7218_/B sky130_fd_sc_hd__xnor2_1
X_4425_ _7539_/B vssd1 vssd1 vccd1 vccd1 _7538_/B sky130_fd_sc_hd__buf_2
X_8193_ _7792_/B _8193_/B vssd1 vssd1 vccd1 vccd1 _8196_/A sky130_fd_sc_hd__and2b_1
X_7144_ _7137_/X _7141_/X _7142_/Y _7143_/X vssd1 vssd1 vccd1 vccd1 _7146_/B sky130_fd_sc_hd__o211ai_1
X_4356_ _4357_/A vssd1 vssd1 vccd1 vccd1 _4356_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4287_ _4289_/A vssd1 vssd1 vccd1 vccd1 _4287_/Y sky130_fd_sc_hd__inv_2
X_7075_ _7075_/A _7075_/B vssd1 vssd1 vccd1 vccd1 _7131_/B sky130_fd_sc_hd__nor2_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6026_ _6026_/A _6151_/S vssd1 vssd1 vccd1 vccd1 _6027_/B sky130_fd_sc_hd__xnor2_1
XFILLER_39_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7977_ _8039_/A _7977_/B vssd1 vssd1 vccd1 vccd1 _7995_/A sky130_fd_sc_hd__xnor2_1
X_6928_ _6917_/X _6921_/B _6918_/A vssd1 vssd1 vccd1 vccd1 _6949_/A sky130_fd_sc_hd__a21o_1
XFILLER_54_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6859_ _6859_/A _7306_/A vssd1 vssd1 vccd1 vccd1 _7289_/B sky130_fd_sc_hd__xnor2_2
XFILLER_22_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8529_ input3/X _8529_/D vssd1 vssd1 vccd1 vccd1 _8529_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8662__78 vssd1 vssd1 vccd1 vccd1 _8662__78/HI _8771_/A sky130_fd_sc_hd__conb_1
XINSDIODE2_71 _8783_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_60 _8776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_82 _8506_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5190_ _8419_/A vssd1 vssd1 vccd1 vccd1 _6426_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_95_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7900_ _7855_/A _7854_/B _7899_/X vssd1 vssd1 vccd1 vccd1 _7901_/B sky130_fd_sc_hd__o21ai_4
XFILLER_48_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7831_ _7826_/Y _7827_/X _7830_/Y _7983_/A vssd1 vssd1 vccd1 vccd1 _7832_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4974_ _4974_/A _4974_/B vssd1 vssd1 vccd1 vccd1 _4974_/X sky130_fd_sc_hd__or2_1
X_7762_ _7803_/A _7921_/B vssd1 vssd1 vccd1 vccd1 _8097_/A sky130_fd_sc_hd__nand2_1
X_6713_ _7248_/B _6781_/A vssd1 vssd1 vccd1 vccd1 _7116_/A sky130_fd_sc_hd__nand2_2
X_7693_ _7693_/A _7798_/B vssd1 vssd1 vccd1 vccd1 _8205_/A sky130_fd_sc_hd__xnor2_2
X_6644_ _7175_/B _6643_/D _6916_/A vssd1 vssd1 vccd1 vccd1 _6896_/C sky130_fd_sc_hd__o21ai_2
XFILLER_32_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6575_ _6575_/A _6575_/B _6575_/C vssd1 vssd1 vccd1 vccd1 _6683_/A sky130_fd_sc_hd__and3_1
X_5526_ _5526_/A _5526_/B vssd1 vssd1 vccd1 vccd1 _5703_/A sky130_fd_sc_hd__nand2_2
X_8314_ _8257_/A _8256_/B _8254_/X vssd1 vssd1 vccd1 vccd1 _8315_/B sky130_fd_sc_hd__a21oi_1
X_8245_ _8245_/A _8245_/B vssd1 vssd1 vccd1 vccd1 _8287_/A sky130_fd_sc_hd__xnor2_1
X_5457_ _5767_/A vssd1 vssd1 vccd1 vccd1 _5828_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4408_ _4408_/A vssd1 vssd1 vccd1 vccd1 _8726_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_59_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8176_ _8176_/A _8176_/B vssd1 vssd1 vccd1 vccd1 _8176_/Y sky130_fd_sc_hd__nor2_1
X_5388_ _5386_/X _5388_/B vssd1 vssd1 vccd1 vccd1 _5563_/B sky130_fd_sc_hd__and2b_2
X_7127_ _7127_/A _7127_/B vssd1 vssd1 vccd1 vccd1 _7151_/B sky130_fd_sc_hd__nor2_2
XFILLER_59_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4339_ _4339_/A vssd1 vssd1 vccd1 vccd1 _4339_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7058_ _7058_/A _7131_/A vssd1 vssd1 vccd1 vccd1 _7077_/B sky130_fd_sc_hd__xnor2_1
XFILLER_75_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6009_ _6010_/A _6010_/B vssd1 vssd1 vccd1 vccd1 _6011_/A sky130_fd_sc_hd__nand2_1
XFILLER_27_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4690_ _7501_/B _4690_/B vssd1 vssd1 vccd1 vccd1 _4691_/C sky130_fd_sc_hd__nand2_1
X_6360_ _6362_/B _6362_/C _6326_/B vssd1 vssd1 vccd1 vccd1 _6360_/Y sky130_fd_sc_hd__o21ai_1
X_5311_ _5311_/A vssd1 vssd1 vccd1 vccd1 _8507_/D sky130_fd_sc_hd__clkinv_2
X_6291_ _6289_/C _6298_/S vssd1 vssd1 vccd1 vccd1 _6295_/A sky130_fd_sc_hd__and2b_1
X_8030_ _8091_/A _8091_/B vssd1 vssd1 vccd1 vccd1 _8031_/B sky130_fd_sc_hd__xor2_1
X_5242_ _8489_/Q _5240_/B _5241_/X vssd1 vssd1 vccd1 vccd1 _5243_/B sky130_fd_sc_hd__o21ai_1
X_5173_ _5173_/A _5173_/B vssd1 vssd1 vccd1 vccd1 _5173_/X sky130_fd_sc_hd__or2_1
Xinput1 active vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_4
XFILLER_68_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7814_ _7926_/A _7983_/A vssd1 vssd1 vccd1 vccd1 _7815_/B sky130_fd_sc_hd__nor2_1
XFILLER_51_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4957_ _5074_/A _5031_/C _4957_/C _4957_/D vssd1 vssd1 vccd1 vccd1 _4957_/X sky130_fd_sc_hd__or4_1
XFILLER_51_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7745_ _7747_/A _7746_/A vssd1 vssd1 vccd1 vccd1 _7866_/A sky130_fd_sc_hd__or2_1
X_4888_ _4969_/A _4955_/B _4884_/X _4887_/X vssd1 vssd1 vccd1 vccd1 _4891_/C sky130_fd_sc_hd__o31a_1
X_7676_ _7796_/B _7676_/B vssd1 vssd1 vccd1 vccd1 _7693_/A sky130_fd_sc_hd__or2_1
X_6627_ _6627_/A _6627_/B _6627_/C vssd1 vssd1 vccd1 vccd1 _6969_/B sky130_fd_sc_hd__nand3_1
X_6558_ _6558_/A _6941_/A vssd1 vssd1 vccd1 vccd1 _6647_/B sky130_fd_sc_hd__and2_1
XFILLER_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6489_ _8550_/Q _8467_/Q vssd1 vssd1 vccd1 vccd1 _6584_/A sky130_fd_sc_hd__xnor2_2
X_5509_ _5509_/A vssd1 vssd1 vccd1 vccd1 _5949_/A sky130_fd_sc_hd__clkbuf_2
X_8228_ _8125_/A _8125_/B _8227_/Y vssd1 vssd1 vccd1 vccd1 _8302_/A sky130_fd_sc_hd__a21bo_1
XFILLER_86_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8159_ _8159_/A _8159_/B vssd1 vssd1 vccd1 vccd1 _8282_/A sky130_fd_sc_hd__xnor2_1
XFILLER_59_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8632__48 vssd1 vssd1 vccd1 vccd1 _8632__48/HI _8741_/A sky130_fd_sc_hd__conb_1
XFILLER_74_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5860_ _5860_/A _5860_/B vssd1 vssd1 vccd1 vccd1 _5860_/Y sky130_fd_sc_hd__nand2_1
XFILLER_18_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4811_ _4811_/A vssd1 vssd1 vccd1 vccd1 _4953_/A sky130_fd_sc_hd__inv_2
XFILLER_21_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5791_ _5978_/A _5855_/B vssd1 vssd1 vccd1 vccd1 _5792_/A sky130_fd_sc_hd__or2_1
XFILLER_33_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4742_ _4755_/A _4742_/B _4765_/A vssd1 vssd1 vccd1 vccd1 _4796_/B sky130_fd_sc_hd__nand3b_2
X_7530_ _7530_/A _7682_/A vssd1 vssd1 vccd1 vccd1 _7530_/Y sky130_fd_sc_hd__nand2_1
X_4673_ _8410_/A _4673_/B vssd1 vssd1 vccd1 vccd1 _8466_/D sky130_fd_sc_hd__nor2_1
X_7461_ _7461_/A _7461_/B vssd1 vssd1 vccd1 vccd1 _7461_/Y sky130_fd_sc_hd__xnor2_1
X_6412_ _6402_/Y _6411_/X _8410_/A vssd1 vssd1 vccd1 vccd1 _8548_/D sky130_fd_sc_hd__a21oi_1
X_7392_ _7388_/A _7388_/B _7386_/A vssd1 vssd1 vccd1 vccd1 _7393_/B sky130_fd_sc_hd__a21oi_1
X_6343_ _8531_/Q _8532_/Q _6343_/C vssd1 vssd1 vccd1 vccd1 _6351_/C sky130_fd_sc_hd__and3_1
X_6274_ _6281_/B _6274_/B vssd1 vssd1 vccd1 vccd1 _6276_/A sky130_fd_sc_hd__and2b_1
X_5225_ _8499_/Q _5224_/X _8501_/Q _8500_/Q vssd1 vssd1 vccd1 vccd1 _5226_/C sky130_fd_sc_hd__o211a_1
X_8013_ _8013_/A _8013_/B vssd1 vssd1 vccd1 vccd1 _8016_/B sky130_fd_sc_hd__xor2_1
XFILLER_96_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5156_ _5156_/A _5156_/B _5156_/C _5156_/D vssd1 vssd1 vccd1 vccd1 _5156_/X sky130_fd_sc_hd__or4_1
X_5087_ _5087_/A _5087_/B vssd1 vssd1 vccd1 vccd1 _5088_/C sky130_fd_sc_hd__or2_1
XFILLER_84_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8777_ _8777_/A _4371_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[24] sky130_fd_sc_hd__ebufn_8
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5989_ _5990_/A _5990_/B _5990_/C vssd1 vssd1 vccd1 vccd1 _5989_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_24_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7728_ _7728_/A _7841_/B _7728_/C vssd1 vssd1 vccd1 vccd1 _7736_/A sky130_fd_sc_hd__and3_1
XFILLER_20_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7659_ _7546_/A _7526_/B _7658_/X vssd1 vssd1 vccd1 vccd1 _7660_/B sky130_fd_sc_hd__o21a_1
XFILLER_79_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5010_ _5010_/A _5169_/A _5010_/C vssd1 vssd1 vccd1 vccd1 _5093_/C sky130_fd_sc_hd__or3_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6961_ _6961_/A _6961_/B vssd1 vssd1 vccd1 vccd1 _6962_/B sky130_fd_sc_hd__and2_1
X_8700_ _8700_/A _4280_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[17] sky130_fd_sc_hd__ebufn_8
XFILLER_19_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6892_ _6892_/A _6990_/A vssd1 vssd1 vccd1 vccd1 _6913_/B sky130_fd_sc_hd__xor2_1
X_5912_ _5994_/A _5912_/B vssd1 vssd1 vccd1 vccd1 _5965_/B sky130_fd_sc_hd__and2_1
XFILLER_34_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5843_ _5843_/A _5843_/B vssd1 vssd1 vccd1 vccd1 _5844_/B sky130_fd_sc_hd__xor2_1
X_8562_ input3/X _8562_/D vssd1 vssd1 vccd1 vccd1 _8562_/Q sky130_fd_sc_hd__dfxtp_1
X_5774_ _5774_/A _5838_/A vssd1 vssd1 vccd1 vccd1 _5826_/A sky130_fd_sc_hd__nor2_2
X_7513_ _7537_/A _7524_/B vssd1 vssd1 vccd1 vccd1 _7768_/A sky130_fd_sc_hd__xnor2_2
X_4725_ _4725_/A _4748_/B _4766_/B _4718_/A vssd1 vssd1 vccd1 vccd1 _4800_/A sky130_fd_sc_hd__or4b_4
X_8493_ input3/X _8493_/D vssd1 vssd1 vccd1 vccd1 _8493_/Q sky130_fd_sc_hd__dfxtp_1
X_4656_ _4659_/A _4655_/X _4656_/S vssd1 vssd1 vccd1 vccd1 _4657_/C sky130_fd_sc_hd__mux2_1
X_7444_ _7518_/A _7417_/A _7443_/Y _7481_/B vssd1 vssd1 vccd1 vccd1 _7444_/X sky130_fd_sc_hd__a31o_1
X_7375_ _6472_/X _8560_/Q _7362_/X _7374_/Y vssd1 vssd1 vccd1 vccd1 _8560_/D sky130_fd_sc_hd__o22a_1
X_4587_ _4748_/B vssd1 vssd1 vccd1 vccd1 _4735_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6326_ _8527_/Q _6326_/B vssd1 vssd1 vccd1 vccd1 _6327_/A sky130_fd_sc_hd__and2b_1
XFILLER_1_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6257_ _6251_/X _6256_/X _4668_/X _8517_/Q vssd1 vssd1 vccd1 vccd1 _8517_/D sky130_fd_sc_hd__o2bb2a_1
X_5208_ _8481_/Q _5217_/B vssd1 vssd1 vccd1 vccd1 _5208_/X sky130_fd_sc_hd__or2_1
X_6188_ _6188_/A _6188_/B vssd1 vssd1 vccd1 vccd1 _6188_/Y sky130_fd_sc_hd__nand2_1
XFILLER_96_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5139_ _5179_/B _4859_/X _5135_/X _4619_/A _5138_/X vssd1 vssd1 vccd1 vccd1 _5139_/X
+ sky130_fd_sc_hd__o221a_1
X_8602__18 vssd1 vssd1 vccd1 vccd1 _8602__18/HI _8697_/A sky130_fd_sc_hd__conb_1
XFILLER_84_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5490_ _5625_/A _5490_/B vssd1 vssd1 vccd1 vccd1 _5604_/B sky130_fd_sc_hd__xor2_1
X_4510_ _4510_/A _5368_/B vssd1 vssd1 vccd1 vccd1 _4511_/B sky130_fd_sc_hd__nand2_1
X_4441_ _7538_/B _4464_/B _4438_/Y _7766_/B vssd1 vssd1 vccd1 vccd1 _4470_/A sky130_fd_sc_hd__o31a_1
XFILLER_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7160_ _7173_/A _7173_/B _7159_/X vssd1 vssd1 vccd1 vccd1 _7162_/A sky130_fd_sc_hd__a21oi_1
X_8668__84 vssd1 vssd1 vccd1 vccd1 _8668__84/HI _8777_/A sky130_fd_sc_hd__conb_1
X_4372_ _4375_/A vssd1 vssd1 vccd1 vccd1 _4372_/Y sky130_fd_sc_hd__inv_2
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6111_ _6111_/A _6111_/B vssd1 vssd1 vccd1 vccd1 _6112_/B sky130_fd_sc_hd__nor2_1
X_7091_ _7143_/A _7088_/Y _7089_/Y _7090_/X vssd1 vssd1 vccd1 vccd1 _7098_/B sky130_fd_sc_hd__o211a_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6042_ _6042_/A _6042_/B _6042_/C vssd1 vssd1 vccd1 vccd1 _6043_/B sky130_fd_sc_hd__nor3_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7993_ _7993_/A _7993_/B vssd1 vssd1 vccd1 vccd1 _7994_/B sky130_fd_sc_hd__nand2_1
X_6944_ _6937_/A _6937_/C _6937_/B vssd1 vssd1 vccd1 vccd1 _6945_/C sky130_fd_sc_hd__a21o_1
XFILLER_54_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6875_ _6875_/A _6875_/B vssd1 vssd1 vccd1 vccd1 _6894_/B sky130_fd_sc_hd__xor2_2
X_5826_ _5826_/A _5840_/B vssd1 vssd1 vccd1 vccd1 _5827_/B sky130_fd_sc_hd__xnor2_2
X_8545_ input3/X _8545_/D vssd1 vssd1 vccd1 vccd1 _8545_/Q sky130_fd_sc_hd__dfxtp_1
X_5757_ _5758_/A _5758_/B vssd1 vssd1 vccd1 vccd1 _5757_/X sky130_fd_sc_hd__or2_1
X_8476_ input3/X _8476_/D vssd1 vssd1 vccd1 vccd1 _8476_/Q sky130_fd_sc_hd__dfxtp_1
X_4708_ _5526_/B _5192_/B _4707_/Y _4663_/B vssd1 vssd1 vccd1 vccd1 _4709_/B sky130_fd_sc_hd__o2bb2a_1
X_5688_ _5793_/A vssd1 vssd1 vccd1 vccd1 _6118_/A sky130_fd_sc_hd__buf_2
X_7427_ _8397_/B _8391_/A _8581_/Q _7426_/Y vssd1 vssd1 vccd1 vccd1 _7427_/X sky130_fd_sc_hd__a31o_1
X_4639_ _4639_/A _4639_/B vssd1 vssd1 vccd1 vccd1 _5046_/A sky130_fd_sc_hd__or2_2
XFILLER_89_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7358_ _7358_/A _7358_/B vssd1 vssd1 vccd1 vccd1 _7359_/B sky130_fd_sc_hd__nand2_1
XFILLER_89_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6309_ _8537_/Q _8536_/Q _8538_/Q vssd1 vssd1 vccd1 vccd1 _6309_/X sky130_fd_sc_hd__a21o_1
X_7289_ _6860_/A _7289_/B vssd1 vssd1 vccd1 vccd1 _7289_/X sky130_fd_sc_hd__and2b_1
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4990_ _5031_/B _5050_/C vssd1 vssd1 vccd1 vccd1 _5018_/C sky130_fd_sc_hd__or2_1
XFILLER_63_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6660_ _6660_/A _6660_/B vssd1 vssd1 vccd1 vccd1 _6661_/B sky130_fd_sc_hd__or2_1
X_6591_ _6591_/A _6591_/B vssd1 vssd1 vccd1 vccd1 _6592_/B sky130_fd_sc_hd__nor2_1
X_5611_ _5610_/B _5722_/A _5628_/A vssd1 vssd1 vccd1 vccd1 _5612_/C sky130_fd_sc_hd__a21bo_1
X_8330_ _8325_/X _8326_/X _8329_/Y vssd1 vssd1 vccd1 vccd1 _8331_/B sky130_fd_sc_hd__a21oi_1
X_5542_ _5426_/A _5406_/B _5541_/X vssd1 vssd1 vccd1 vccd1 _5543_/B sky130_fd_sc_hd__o21a_1
X_8261_ _7607_/Y _8063_/B _8260_/X vssd1 vssd1 vccd1 vccd1 _8263_/A sky130_fd_sc_hd__o21a_1
X_5473_ _5560_/A _5560_/B vssd1 vssd1 vccd1 vccd1 _5561_/A sky130_fd_sc_hd__nor2_1
X_7212_ _7212_/A _7212_/B vssd1 vssd1 vccd1 vccd1 _7213_/B sky130_fd_sc_hd__xor2_1
X_4424_ _8472_/Q vssd1 vssd1 vccd1 vccd1 _7539_/B sky130_fd_sc_hd__inv_2
X_8192_ _8202_/A _8192_/B vssd1 vssd1 vccd1 vccd1 _8192_/X sky130_fd_sc_hd__xor2_1
X_7143_ _7143_/A _7143_/B _7143_/C vssd1 vssd1 vccd1 vccd1 _7143_/X sky130_fd_sc_hd__or3_1
X_4355_ _4357_/A vssd1 vssd1 vccd1 vccd1 _4355_/Y sky130_fd_sc_hd__inv_2
X_7074_ _7116_/B _7126_/B _7008_/B _7126_/A vssd1 vssd1 vccd1 vccd1 _7075_/B sky130_fd_sc_hd__o211a_1
XFILLER_58_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4286_ _4289_/A vssd1 vssd1 vccd1 vccd1 _4286_/Y sky130_fd_sc_hd__inv_2
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6025_ _6025_/A _6025_/B vssd1 vssd1 vccd1 vccd1 _6151_/S sky130_fd_sc_hd__nor2_2
XFILLER_73_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7976_ _7976_/A _7976_/B vssd1 vssd1 vccd1 vccd1 _7977_/B sky130_fd_sc_hd__xor2_2
XFILLER_81_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6927_ _6990_/A _6990_/B vssd1 vssd1 vccd1 vccd1 _6991_/A sky130_fd_sc_hd__nand2_2
X_6858_ _6858_/A _6858_/B vssd1 vssd1 vccd1 vccd1 _7306_/A sky130_fd_sc_hd__and2_1
XFILLER_50_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5809_ _5809_/A _5809_/B _5809_/C vssd1 vssd1 vccd1 vccd1 _5810_/B sky130_fd_sc_hd__nand3_1
X_6789_ _7321_/A _7321_/B vssd1 vssd1 vccd1 vccd1 _6789_/Y sky130_fd_sc_hd__xnor2_1
X_8528_ input3/X _8528_/D vssd1 vssd1 vccd1 vccd1 _8528_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8459_ input3/X _8459_/D vssd1 vssd1 vccd1 vccd1 _8459_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_61 _8776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_50 _8767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_72 _8784_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_83 _8506_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8638__54 vssd1 vssd1 vccd1 vccd1 _8638__54/HI _8747_/A sky130_fd_sc_hd__conb_1
XFILLER_95_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7830_ _7926_/A _7830_/B vssd1 vssd1 vccd1 vccd1 _7830_/Y sky130_fd_sc_hd__nor2_1
XFILLER_36_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4973_ _4973_/A _5147_/A _5020_/C _5058_/B vssd1 vssd1 vccd1 vccd1 _4974_/B sky130_fd_sc_hd__or4_1
XFILLER_63_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7761_ _7822_/B vssd1 vssd1 vccd1 vccd1 _7921_/B sky130_fd_sc_hd__clkbuf_2
X_6712_ _6939_/B _7323_/B vssd1 vssd1 vccd1 vccd1 _6781_/A sky130_fd_sc_hd__nor2_2
X_7692_ _7679_/A _8023_/A _7694_/B _7691_/A vssd1 vssd1 vccd1 vccd1 _7798_/B sky130_fd_sc_hd__a31o_1
X_6643_ _6977_/A _6829_/A _6643_/C _6643_/D vssd1 vssd1 vccd1 vccd1 _6916_/A sky130_fd_sc_hd__nand4_2
X_6574_ _6521_/X _6574_/B vssd1 vssd1 vccd1 vccd1 _6575_/A sky130_fd_sc_hd__and2b_1
X_8313_ _8245_/A _8245_/B _8312_/X vssd1 vssd1 vccd1 vccd1 _8315_/A sky130_fd_sc_hd__a21oi_1
X_5525_ _5978_/A _5855_/A vssd1 vssd1 vccd1 vccd1 _5541_/B sky130_fd_sc_hd__nor2_1
X_8244_ _8244_/A vssd1 vssd1 vccd1 vccd1 _8245_/B sky130_fd_sc_hd__inv_2
X_5456_ _5607_/A vssd1 vssd1 vccd1 vccd1 _5767_/A sky130_fd_sc_hd__clkbuf_2
X_4407_ _4469_/A _4642_/A vssd1 vssd1 vccd1 vccd1 _4408_/A sky130_fd_sc_hd__or2_1
X_5387_ _8470_/Q _8512_/Q vssd1 vssd1 vccd1 vccd1 _5388_/B sky130_fd_sc_hd__or2b_1
X_8175_ _8292_/A _8359_/B vssd1 vssd1 vccd1 vccd1 _8364_/A sky130_fd_sc_hd__xnor2_1
X_7126_ _7126_/A _7126_/B _7126_/C _7126_/D vssd1 vssd1 vccd1 vccd1 _7127_/B sky130_fd_sc_hd__and4_1
X_4338_ _4339_/A vssd1 vssd1 vccd1 vccd1 _4338_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4269_ _4270_/A vssd1 vssd1 vccd1 vccd1 _4269_/Y sky130_fd_sc_hd__inv_2
X_7057_ _7057_/A _7057_/B vssd1 vssd1 vccd1 vccd1 _7077_/A sky130_fd_sc_hd__nand2_1
XFILLER_55_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6008_ _6008_/A _6008_/B vssd1 vssd1 vccd1 vccd1 _6010_/B sky130_fd_sc_hd__xor2_1
XFILLER_27_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7959_ _7959_/A _7958_/X vssd1 vssd1 vccd1 vccd1 _7967_/A sky130_fd_sc_hd__or2b_1
XFILLER_27_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6290_ _5333_/A _6288_/Y _6298_/S _5332_/A _6286_/B vssd1 vssd1 vccd1 vccd1 _8524_/D
+ sky130_fd_sc_hd__a32o_1
X_5310_ _6293_/A _6286_/B _5306_/X _5309_/Y _4510_/A vssd1 vssd1 vccd1 vccd1 _5311_/A
+ sky130_fd_sc_hd__o311a_1
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5241_ _5260_/A vssd1 vssd1 vccd1 vccd1 _5241_/X sky130_fd_sc_hd__buf_2
X_5172_ _4909_/B _5151_/C _5169_/X _5171_/X vssd1 vssd1 vccd1 vccd1 _5173_/B sky130_fd_sc_hd__o31a_1
XFILLER_96_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput2 io_in[10] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__clkbuf_2
XFILLER_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7813_ _7813_/A vssd1 vssd1 vccd1 vccd1 _7926_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_24_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7744_ _7744_/A _7744_/B vssd1 vssd1 vccd1 vccd1 _7750_/B sky130_fd_sc_hd__nand2_1
X_4956_ _5101_/S _5151_/B _4956_/C _5132_/D vssd1 vssd1 vccd1 vccd1 _4957_/D sky130_fd_sc_hd__or4_1
X_4887_ _5101_/S _5012_/C _4887_/C vssd1 vssd1 vccd1 vccd1 _4887_/X sky130_fd_sc_hd__or3_1
X_7675_ _7796_/A _7674_/C _7674_/A vssd1 vssd1 vccd1 vccd1 _7676_/B sky130_fd_sc_hd__o21a_1
X_6626_ _6914_/B _6977_/A _6844_/S vssd1 vssd1 vccd1 vccd1 _6626_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_20_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6557_ _6557_/A vssd1 vssd1 vccd1 vccd1 _6941_/A sky130_fd_sc_hd__clkbuf_4
X_5508_ _5609_/C _5825_/B _5825_/C vssd1 vssd1 vccd1 vccd1 _5509_/A sky130_fd_sc_hd__or3_1
X_6488_ _8551_/Q _8468_/Q vssd1 vssd1 vccd1 vccd1 _6501_/B sky130_fd_sc_hd__xnor2_2
XFILLER_10_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5439_ _8458_/Q vssd1 vssd1 vccd1 vccd1 _7559_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_10_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8227_ _8227_/A _8348_/A vssd1 vssd1 vccd1 vccd1 _8227_/Y sky130_fd_sc_hd__nand2_1
XFILLER_87_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8158_ _8277_/B _8270_/A vssd1 vssd1 vccd1 vccd1 _8159_/B sky130_fd_sc_hd__xnor2_1
XFILLER_87_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7109_ _7109_/A _7109_/B vssd1 vssd1 vccd1 vccd1 _7129_/B sky130_fd_sc_hd__xnor2_1
XFILLER_74_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8089_ _8080_/A _8080_/B _8088_/Y vssd1 vssd1 vccd1 vccd1 _8218_/B sky130_fd_sc_hd__a21o_1
XFILLER_47_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8608__24 vssd1 vssd1 vccd1 vccd1 _8608__24/HI _8703_/A sky130_fd_sc_hd__conb_1
XFILLER_78_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4810_ _5112_/A _4969_/A vssd1 vssd1 vccd1 vccd1 _4985_/A sky130_fd_sc_hd__or2_1
XFILLER_33_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5790_ _5581_/A _6183_/S _5708_/X vssd1 vssd1 vccd1 vccd1 _5794_/A sky130_fd_sc_hd__o21a_1
X_4741_ _5144_/B _4741_/B vssd1 vssd1 vccd1 vccd1 _4765_/A sky130_fd_sc_hd__or2_2
XFILLER_14_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4672_ _4670_/A _5192_/B _4671_/X vssd1 vssd1 vccd1 vccd1 _4673_/B sky130_fd_sc_hd__a21oi_1
X_7460_ _7494_/A _7454_/B _7453_/A vssd1 vssd1 vccd1 vccd1 _7461_/B sky130_fd_sc_hd__o21a_1
X_6411_ _6407_/X _6409_/X _7403_/A _8565_/Q vssd1 vssd1 vccd1 vccd1 _6411_/X sky130_fd_sc_hd__a211o_1
X_7391_ _7391_/A _7391_/B vssd1 vssd1 vccd1 vccd1 _7393_/A sky130_fd_sc_hd__nand2_1
X_6342_ _6319_/D _6343_/C _6341_/Y vssd1 vssd1 vccd1 vccd1 _8531_/D sky130_fd_sc_hd__a21oi_1
X_6273_ _6270_/A _5332_/X _5333_/X _6272_/Y vssd1 vssd1 vccd1 vccd1 _8521_/D sky130_fd_sc_hd__a22o_1
X_5224_ _8497_/Q _8496_/Q _5223_/X _8498_/Q vssd1 vssd1 vccd1 vccd1 _5224_/X sky130_fd_sc_hd__a31o_1
X_8012_ _8012_/A _8012_/B vssd1 vssd1 vccd1 vccd1 _8013_/B sky130_fd_sc_hd__xor2_1
X_5155_ _5164_/B _4868_/X _5148_/C _4937_/X _4989_/A vssd1 vssd1 vccd1 vccd1 _5156_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_69_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5086_ _5009_/C _5085_/X _4848_/A vssd1 vssd1 vccd1 vccd1 _5089_/C sky130_fd_sc_hd__o21a_1
XFILLER_56_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8776_ _8776_/A _4369_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[23] sky130_fd_sc_hd__ebufn_8
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5988_ _6115_/B _5988_/B vssd1 vssd1 vccd1 vccd1 _5990_/C sky130_fd_sc_hd__xor2_1
XFILLER_24_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4939_ _5053_/B _4939_/B vssd1 vssd1 vccd1 vccd1 _4939_/X sky130_fd_sc_hd__or2_1
X_7727_ _7726_/B _7841_/A _7747_/A vssd1 vssd1 vccd1 vccd1 _7728_/C sky130_fd_sc_hd__a21bo_1
XFILLER_20_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7658_ _7921_/A _7658_/B vssd1 vssd1 vccd1 vccd1 _7658_/X sky130_fd_sc_hd__or2_1
X_6609_ _6609_/A _6609_/B _6609_/C vssd1 vssd1 vccd1 vccd1 _6640_/A sky130_fd_sc_hd__and3_1
XFILLER_21_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7589_ _7844_/A vssd1 vssd1 vccd1 vccd1 _8317_/B sky130_fd_sc_hd__buf_2
XFILLER_87_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6960_ _6961_/A _6960_/B _6960_/C vssd1 vssd1 vccd1 vccd1 _6961_/B sky130_fd_sc_hd__nand3_1
XFILLER_66_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5911_ _5911_/A _5911_/B vssd1 vssd1 vccd1 vccd1 _5912_/B sky130_fd_sc_hd__or2_1
X_6891_ _6891_/A _6891_/B vssd1 vssd1 vccd1 vccd1 _7280_/B sky130_fd_sc_hd__xnor2_1
X_5842_ _5927_/A _5842_/B vssd1 vssd1 vccd1 vccd1 _5843_/B sky130_fd_sc_hd__xnor2_1
XFILLER_34_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8561_ input3/X _8561_/D vssd1 vssd1 vccd1 vccd1 _8561_/Q sky130_fd_sc_hd__dfxtp_2
X_5773_ _5821_/A _5821_/B vssd1 vssd1 vccd1 vccd1 _5782_/A sky130_fd_sc_hd__xnor2_4
X_4724_ _4882_/A _4796_/A _4899_/B vssd1 vssd1 vccd1 vccd1 _4782_/B sky130_fd_sc_hd__o21a_1
X_7512_ _7805_/A vssd1 vssd1 vccd1 vccd1 _7804_/A sky130_fd_sc_hd__clkbuf_2
X_8492_ input3/X _8492_/D vssd1 vssd1 vccd1 vccd1 _8492_/Q sky130_fd_sc_hd__dfxtp_1
X_4655_ _4655_/A _5180_/A vssd1 vssd1 vccd1 vccd1 _4655_/X sky130_fd_sc_hd__or2b_1
X_7443_ _7501_/A _7452_/A _8573_/Q vssd1 vssd1 vccd1 vccd1 _7443_/Y sky130_fd_sc_hd__o21ai_1
X_7374_ _7372_/X _7373_/Y _7366_/B vssd1 vssd1 vccd1 vccd1 _7374_/Y sky130_fd_sc_hd__a21boi_1
X_4586_ _8465_/Q vssd1 vssd1 vccd1 vccd1 _4748_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6325_ _6389_/B vssd1 vssd1 vccd1 vccd1 _6326_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_88_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6256_ _6264_/A _6264_/B _6264_/C _6256_/D vssd1 vssd1 vccd1 vccd1 _6256_/X sky130_fd_sc_hd__or4_1
X_5207_ _5207_/A vssd1 vssd1 vccd1 vccd1 _5217_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6187_ _6146_/A _6146_/B _6144_/A vssd1 vssd1 vccd1 vccd1 _6192_/A sky130_fd_sc_hd__o21ai_1
X_8599__15 vssd1 vssd1 vccd1 vccd1 _8599__15/HI _8694_/A sky130_fd_sc_hd__conb_1
XFILLER_96_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5138_ _5138_/A _5138_/B _5138_/C _5138_/D vssd1 vssd1 vccd1 vccd1 _5138_/X sky130_fd_sc_hd__or4_1
XFILLER_57_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5069_ _5069_/A _5179_/A _5132_/A _5136_/C vssd1 vssd1 vccd1 vccd1 _5069_/X sky130_fd_sc_hd__or4_1
XFILLER_72_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8759_ _8759_/A _4339_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[6] sky130_fd_sc_hd__ebufn_8
XFILLER_12_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4440_ _7644_/B vssd1 vssd1 vccd1 vccd1 _7766_/B sky130_fd_sc_hd__clkbuf_4
X_4371_ _4375_/A vssd1 vssd1 vccd1 vccd1 _4371_/Y sky130_fd_sc_hd__inv_2
X_6110_ _6110_/A _6110_/B _6110_/C vssd1 vssd1 vccd1 vccd1 _6111_/B sky130_fd_sc_hd__nor3_1
X_7090_ _7017_/B _7019_/C _7021_/Y _7022_/X vssd1 vssd1 vccd1 vccd1 _7090_/X sky130_fd_sc_hd__a211o_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6041_ _6042_/A _6042_/B _6042_/C vssd1 vssd1 vccd1 vccd1 _6043_/A sky130_fd_sc_hd__o21a_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7992_ _7993_/A _7993_/B vssd1 vssd1 vccd1 vccd1 _7994_/A sky130_fd_sc_hd__or2_1
X_6943_ _7009_/A _7009_/B vssd1 vssd1 vccd1 vccd1 _6945_/B sky130_fd_sc_hd__and2b_1
X_6874_ _6874_/A _6874_/B _6874_/C vssd1 vssd1 vccd1 vccd1 _6880_/A sky130_fd_sc_hd__nand3_1
XFILLER_22_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5825_ _5825_/A _5825_/B _5825_/C vssd1 vssd1 vccd1 vccd1 _5840_/B sky130_fd_sc_hd__or3_2
X_8544_ input3/X _8544_/D vssd1 vssd1 vccd1 vccd1 _8544_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5756_ _5743_/A _5753_/Y _5754_/X _5755_/X vssd1 vssd1 vccd1 vccd1 _5783_/A sky130_fd_sc_hd__a31o_2
X_8475_ input3/X _8475_/D vssd1 vssd1 vccd1 vccd1 _8475_/Q sky130_fd_sc_hd__dfxtp_1
X_4707_ _5526_/B _4707_/B vssd1 vssd1 vccd1 vccd1 _4707_/Y sky130_fd_sc_hd__xnor2_1
X_5687_ _5651_/A _5900_/B _5795_/A vssd1 vssd1 vccd1 vccd1 _5793_/A sky130_fd_sc_hd__mux2_2
X_4638_ _4638_/A _4950_/A vssd1 vssd1 vccd1 vccd1 _4639_/B sky130_fd_sc_hd__nor2_1
X_7426_ _8415_/A vssd1 vssd1 vccd1 vccd1 _7426_/Y sky130_fd_sc_hd__inv_2
X_7357_ _7365_/A _7366_/B vssd1 vssd1 vccd1 vccd1 _7357_/X sky130_fd_sc_hd__and2_1
X_4569_ _4569_/A vssd1 vssd1 vccd1 vccd1 _8450_/D sky130_fd_sc_hd__clkbuf_1
X_6308_ _6351_/A _8532_/Q _6307_/X _8534_/Q vssd1 vssd1 vccd1 vccd1 _6308_/X sky130_fd_sc_hd__a211o_1
X_7288_ _7288_/A _7288_/B vssd1 vssd1 vccd1 vccd1 _7303_/A sky130_fd_sc_hd__xnor2_1
XFILLER_1_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6239_ _6239_/A _6239_/B _6239_/C vssd1 vssd1 vccd1 vccd1 _6239_/X sky130_fd_sc_hd__and3_1
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6590_ _6590_/A _8472_/Q vssd1 vssd1 vccd1 vccd1 _6591_/A sky130_fd_sc_hd__nor2_1
X_5610_ _5628_/A _5610_/B _5722_/A vssd1 vssd1 vccd1 vccd1 _5722_/B sky130_fd_sc_hd__nand3b_1
X_5541_ _5800_/A _5541_/B vssd1 vssd1 vccd1 vccd1 _5541_/X sky130_fd_sc_hd__or2_1
XFILLER_31_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8260_ _8260_/A _8260_/B _8260_/C vssd1 vssd1 vccd1 vccd1 _8260_/X sky130_fd_sc_hd__or3_1
X_7211_ _7211_/A _7211_/B _7211_/C vssd1 vssd1 vccd1 vccd1 _7226_/A sky130_fd_sc_hd__nor3_2
X_5472_ _5472_/A _5472_/B vssd1 vssd1 vccd1 vccd1 _5560_/B sky130_fd_sc_hd__xnor2_1
X_4423_ _4698_/A _4698_/B _4715_/A _4438_/A vssd1 vssd1 vccd1 vccd1 _4706_/B sky130_fd_sc_hd__and4_1
X_8191_ _8292_/A _8191_/B vssd1 vssd1 vccd1 vccd1 _8192_/B sky130_fd_sc_hd__nor2_1
X_7142_ _7143_/A _7143_/C _7143_/B vssd1 vssd1 vccd1 vccd1 _7142_/Y sky130_fd_sc_hd__o21ai_1
X_4354_ _4357_/A vssd1 vssd1 vccd1 vccd1 _4354_/Y sky130_fd_sc_hd__inv_2
X_7073_ _7123_/A _7228_/A vssd1 vssd1 vccd1 vccd1 _7126_/B sky130_fd_sc_hd__or2_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4285_ _4289_/A vssd1 vssd1 vccd1 vccd1 _4285_/Y sky130_fd_sc_hd__inv_2
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6024_ _5949_/A _6150_/A _5778_/X vssd1 vssd1 vccd1 vccd1 _6135_/A sky130_fd_sc_hd__o21a_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7975_ _8046_/A _7975_/B vssd1 vssd1 vccd1 vccd1 _7976_/B sky130_fd_sc_hd__nor2_1
XFILLER_81_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6926_ _6926_/A _6926_/B vssd1 vssd1 vccd1 vccd1 _6990_/B sky130_fd_sc_hd__xnor2_1
XFILLER_81_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6857_ _6857_/A _6857_/B vssd1 vssd1 vccd1 vccd1 _6859_/A sky130_fd_sc_hd__xnor2_1
XFILLER_22_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6788_ _7202_/B _6819_/B _6787_/X vssd1 vssd1 vccd1 vccd1 _7321_/B sky130_fd_sc_hd__o21a_1
X_5808_ _5809_/A _5809_/C _5809_/B vssd1 vssd1 vccd1 vccd1 _5870_/A sky130_fd_sc_hd__a21o_1
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8527_ input3/X _8527_/D vssd1 vssd1 vccd1 vccd1 _8527_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5739_ _5739_/A _5765_/A vssd1 vssd1 vccd1 vccd1 _5740_/B sky130_fd_sc_hd__xnor2_1
XFILLER_13_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8458_ input3/X _8458_/D vssd1 vssd1 vccd1 vccd1 _8458_/Q sky130_fd_sc_hd__dfxtp_1
X_7409_ _7404_/A _7408_/X _7409_/S vssd1 vssd1 vccd1 vccd1 _7410_/C sky130_fd_sc_hd__mux2_1
X_8389_ _8387_/Y _7448_/X _8388_/Y vssd1 vssd1 vccd1 vccd1 _8581_/D sky130_fd_sc_hd__o21a_1
XFILLER_89_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_51 _8767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_40 _8716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_73 _8784_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_84 _4390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_62 _8777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8653__69 vssd1 vssd1 vccd1 vccd1 _8653__69/HI _8762_/A sky130_fd_sc_hd__conb_1
XFILLER_95_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4972_ _4972_/A _5112_/D vssd1 vssd1 vccd1 vccd1 _4974_/A sky130_fd_sc_hd__or2_1
X_7760_ _7783_/A _7783_/B vssd1 vssd1 vccd1 vccd1 _7818_/A sky130_fd_sc_hd__or2_1
X_6711_ _7001_/B _7067_/B vssd1 vssd1 vccd1 vccd1 _6938_/A sky130_fd_sc_hd__nand2_1
X_7691_ _7691_/A _7691_/B vssd1 vssd1 vccd1 vccd1 _7694_/B sky130_fd_sc_hd__nor2_1
X_6642_ _6640_/A _6622_/B _7032_/B vssd1 vssd1 vccd1 vccd1 _6643_/C sky130_fd_sc_hd__o21ai_1
XFILLER_32_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6573_ _6714_/C vssd1 vssd1 vccd1 vccd1 _7323_/B sky130_fd_sc_hd__clkbuf_2
X_8312_ _8242_/B _8312_/B vssd1 vssd1 vccd1 vccd1 _8312_/X sky130_fd_sc_hd__and2b_1
XFILLER_8_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5524_ _5524_/A _5524_/B vssd1 vssd1 vccd1 vccd1 _5978_/A sky130_fd_sc_hd__xnor2_4
X_8243_ _8023_/B _8112_/B _8110_/Y vssd1 vssd1 vccd1 vccd1 _8244_/A sky130_fd_sc_hd__a21oi_1
X_5455_ _5455_/A _5455_/B vssd1 vssd1 vccd1 vccd1 _5607_/A sky130_fd_sc_hd__xnor2_1
X_4406_ _5178_/B _4638_/A _4949_/A vssd1 vssd1 vccd1 vccd1 _4642_/A sky130_fd_sc_hd__and3_1
X_8174_ _8291_/A _8174_/B vssd1 vssd1 vccd1 vccd1 _8359_/B sky130_fd_sc_hd__nand2_1
X_7125_ _7126_/A _7126_/C _7126_/D _7126_/B vssd1 vssd1 vccd1 vccd1 _7127_/A sky130_fd_sc_hd__a22oi_1
X_5386_ _8512_/Q _7506_/B vssd1 vssd1 vccd1 vccd1 _5386_/X sky130_fd_sc_hd__and2b_1
XFILLER_86_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4337_ _4339_/A vssd1 vssd1 vccd1 vccd1 _4337_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4268_ _4270_/A vssd1 vssd1 vccd1 vccd1 _4268_/Y sky130_fd_sc_hd__inv_2
X_7056_ _7109_/A _7109_/B vssd1 vssd1 vccd1 vccd1 _7060_/A sky130_fd_sc_hd__nand2_1
XFILLER_74_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6007_ _6134_/A _6007_/B vssd1 vssd1 vccd1 vccd1 _6008_/B sky130_fd_sc_hd__or2_1
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7958_ _7896_/Y _7893_/B _7956_/X _7945_/B vssd1 vssd1 vccd1 vccd1 _7958_/X sky130_fd_sc_hd__a211o_1
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6909_ _6909_/A _6909_/B _6909_/C vssd1 vssd1 vccd1 vccd1 _6910_/B sky130_fd_sc_hd__or3_1
X_7889_ _7888_/X _7845_/X _7844_/Y _7860_/A vssd1 vssd1 vccd1 vccd1 _7944_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_23_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5240_ _8489_/Q _5240_/B vssd1 vssd1 vccd1 vccd1 _5246_/C sky130_fd_sc_hd__and2_1
XFILLER_5_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5171_ _5171_/A _5171_/B _5171_/C _5171_/D vssd1 vssd1 vccd1 vccd1 _5171_/X sky130_fd_sc_hd__or4_1
XFILLER_96_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput3 wb_clk_i vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_16
XFILLER_64_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7812_ _7932_/A _7932_/B vssd1 vssd1 vccd1 vccd1 _7817_/A sky130_fd_sc_hd__xnor2_1
XFILLER_36_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4955_ _4955_/A _4955_/B _4995_/C _5138_/B vssd1 vssd1 vccd1 vccd1 _4955_/X sky130_fd_sc_hd__or4_1
XFILLER_51_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7743_ _7743_/A _7861_/A vssd1 vssd1 vccd1 vccd1 _7750_/A sky130_fd_sc_hd__or2_1
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4886_ _4886_/A _4993_/B _4886_/C _4886_/D vssd1 vssd1 vccd1 vccd1 _4887_/C sky130_fd_sc_hd__or4_1
X_7674_ _7674_/A _7796_/A _7674_/C vssd1 vssd1 vccd1 vccd1 _7796_/B sky130_fd_sc_hd__nor3_1
X_6625_ _6632_/A _6842_/B vssd1 vssd1 vccd1 vccd1 _6844_/S sky130_fd_sc_hd__nor2_1
X_6556_ _6929_/A vssd1 vssd1 vccd1 vccd1 _6660_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5507_ _5764_/C vssd1 vssd1 vccd1 vccd1 _5825_/C sky130_fd_sc_hd__clkbuf_2
X_6487_ _6506_/A vssd1 vssd1 vccd1 vccd1 _7202_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_8226_ _8104_/A _8224_/Y _8225_/Y vssd1 vssd1 vccd1 vccd1 _8237_/A sky130_fd_sc_hd__o21ai_1
X_5438_ _8457_/Q _8520_/Q vssd1 vssd1 vccd1 vccd1 _5455_/A sky130_fd_sc_hd__or2b_1
XFILLER_87_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5369_ _5368_/B _5368_/C _5526_/A vssd1 vssd1 vccd1 vccd1 _5370_/C sky130_fd_sc_hd__o21ai_1
X_8157_ _8072_/A _8156_/A _8277_/A vssd1 vssd1 vccd1 vccd1 _8270_/A sky130_fd_sc_hd__a21oi_1
X_7108_ _7152_/A _7152_/B vssd1 vssd1 vccd1 vccd1 _7153_/A sky130_fd_sc_hd__or2_1
XFILLER_59_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8088_ _8088_/A _8088_/B vssd1 vssd1 vccd1 vccd1 _8088_/Y sky130_fd_sc_hd__nor2_1
XFILLER_87_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7039_ _7043_/A _7039_/B vssd1 vssd1 vccd1 vccd1 _7102_/A sky130_fd_sc_hd__nor2_2
XFILLER_59_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8623__39 vssd1 vssd1 vccd1 vccd1 _8623__39/HI _8718_/A sky130_fd_sc_hd__conb_1
XFILLER_78_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4740_ _5380_/B _7498_/B _4740_/C vssd1 vssd1 vccd1 vccd1 _4741_/B sky130_fd_sc_hd__and3_1
X_4671_ _4671_/A _4671_/B _4780_/B vssd1 vssd1 vccd1 vccd1 _4671_/X sky130_fd_sc_hd__and3_1
X_6410_ _8566_/Q vssd1 vssd1 vccd1 vccd1 _7403_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7390_ _7390_/A _6562_/B vssd1 vssd1 vccd1 vccd1 _7391_/B sky130_fd_sc_hd__or2b_1
X_6341_ _6319_/D _6343_/C _6326_/B vssd1 vssd1 vccd1 vccd1 _6341_/Y sky130_fd_sc_hd__o21ai_1
X_6272_ _8520_/Q _6272_/B vssd1 vssd1 vccd1 vccd1 _6272_/Y sky130_fd_sc_hd__xnor2_1
X_5223_ _8493_/Q _8492_/Q _5221_/X _6396_/D _8495_/Q vssd1 vssd1 vccd1 vccd1 _5223_/X
+ sky130_fd_sc_hd__a311o_1
X_8011_ _8011_/A _8011_/B vssd1 vssd1 vccd1 vccd1 _8012_/B sky130_fd_sc_hd__nand2_1
X_5154_ _5135_/A _5093_/B _5169_/A _5033_/C _5153_/X vssd1 vssd1 vccd1 vccd1 _5154_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_69_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5085_ _5087_/A _5104_/C _5104_/D vssd1 vssd1 vccd1 vccd1 _5085_/X sky130_fd_sc_hd__or3_1
XFILLER_37_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8775_ _8775_/A _4368_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[22] sky130_fd_sc_hd__ebufn_8
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5987_ _5987_/A _5987_/B vssd1 vssd1 vccd1 vccd1 _5988_/B sky130_fd_sc_hd__xnor2_1
X_4938_ _4938_/A _5030_/C vssd1 vssd1 vccd1 vccd1 _4939_/B sky130_fd_sc_hd__or2_1
X_7726_ _7747_/A _7726_/B _7841_/A vssd1 vssd1 vccd1 vccd1 _7841_/B sky130_fd_sc_hd__nand3b_1
X_4869_ _4969_/B _4869_/B vssd1 vssd1 vccd1 vccd1 _5039_/B sky130_fd_sc_hd__or2_1
X_7657_ _7657_/A vssd1 vssd1 vccd1 vccd1 _7783_/A sky130_fd_sc_hd__clkbuf_2
X_6608_ _7033_/A _6842_/B vssd1 vssd1 vccd1 vccd1 _6804_/A sky130_fd_sc_hd__nor2_2
X_7588_ _7677_/A _7677_/B vssd1 vssd1 vccd1 vccd1 _7678_/A sky130_fd_sc_hd__nor2_1
X_6539_ _6539_/A _6539_/B vssd1 vssd1 vccd1 vccd1 _6609_/A sky130_fd_sc_hd__nor2_1
XFILLER_79_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8209_ _8209_/A _8209_/B vssd1 vssd1 vccd1 vccd1 _8361_/B sky130_fd_sc_hd__xnor2_2
XFILLER_87_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5910_ _5911_/A _5911_/B vssd1 vssd1 vccd1 vccd1 _5994_/A sky130_fd_sc_hd__nand2_1
XFILLER_19_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6890_ _6890_/A _7277_/A vssd1 vssd1 vccd1 vccd1 _6891_/B sky130_fd_sc_hd__xnor2_1
XFILLER_22_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5841_ _5841_/A _5841_/B vssd1 vssd1 vccd1 vccd1 _5842_/B sky130_fd_sc_hd__xor2_2
X_8560_ input3/X _8560_/D vssd1 vssd1 vccd1 vccd1 _8560_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5772_ _6021_/A _5772_/B vssd1 vssd1 vccd1 vccd1 _5821_/B sky130_fd_sc_hd__xnor2_2
X_4723_ _4748_/D _4735_/B _4761_/B _4735_/A vssd1 vssd1 vccd1 vccd1 _4899_/B sky130_fd_sc_hd__or4b_4
X_8491_ input3/X _8491_/D vssd1 vssd1 vccd1 vccd1 _8491_/Q sky130_fd_sc_hd__dfxtp_1
X_7511_ _7824_/A _7546_/A vssd1 vssd1 vccd1 vccd1 _7679_/A sky130_fd_sc_hd__nor2_1
X_7442_ _7539_/A _7438_/Y _7477_/A _7766_/A vssd1 vssd1 vccd1 vccd1 _7442_/Y sky130_fd_sc_hd__a31oi_1
X_4654_ _4652_/X _4653_/Y _4602_/X vssd1 vssd1 vccd1 vccd1 _8462_/D sky130_fd_sc_hd__o21a_1
X_7373_ _7372_/B _7372_/C _7372_/A vssd1 vssd1 vccd1 vccd1 _7373_/Y sky130_fd_sc_hd__o21ai_1
X_4585_ _5135_/A vssd1 vssd1 vccd1 vccd1 _4592_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6324_ _6328_/A _7462_/A vssd1 vssd1 vccd1 vccd1 _6389_/B sky130_fd_sc_hd__and2_1
X_6255_ _6259_/B _6255_/B vssd1 vssd1 vccd1 vccd1 _6256_/D sky130_fd_sc_hd__or2_1
X_5206_ _8579_/Q _5202_/X _5205_/X _5200_/X vssd1 vssd1 vccd1 vccd1 _8480_/D sky130_fd_sc_hd__o211a_1
XFILLER_67_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6186_ _6186_/A _6186_/B vssd1 vssd1 vccd1 vccd1 _6194_/A sky130_fd_sc_hd__xnor2_1
X_5137_ _5132_/B _4987_/A _5136_/X _5059_/X vssd1 vssd1 vccd1 vccd1 _5138_/D sky130_fd_sc_hd__o31a_1
X_5068_ _4863_/X _5062_/X _5067_/X _5109_/A vssd1 vssd1 vccd1 vccd1 _5068_/X sky130_fd_sc_hd__o211a_1
XFILLER_29_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8758_ _8758_/A _4341_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[5] sky130_fd_sc_hd__ebufn_8
XFILLER_40_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7709_ _7709_/A vssd1 vssd1 vccd1 vccd1 _8381_/A sky130_fd_sc_hd__inv_2
XFILLER_12_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8689_ _8689_/A _4266_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[6] sky130_fd_sc_hd__ebufn_8
XFILLER_32_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4370_ _4382_/A vssd1 vssd1 vccd1 vccd1 _4375_/A sky130_fd_sc_hd__buf_2
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6040_ _6040_/A _6040_/B vssd1 vssd1 vccd1 vccd1 _6042_/C sky130_fd_sc_hd__xnor2_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7991_ _7991_/A _7991_/B vssd1 vssd1 vccd1 vccd1 _7993_/B sky130_fd_sc_hd__xnor2_1
XFILLER_81_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6942_ _7202_/B _7055_/A _6786_/B vssd1 vssd1 vccd1 vccd1 _7009_/B sky130_fd_sc_hd__a21oi_2
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6873_ _6873_/A _6873_/B vssd1 vssd1 vccd1 vccd1 _6890_/A sky130_fd_sc_hd__xor2_2
X_5824_ _5824_/A _5824_/B _5824_/C vssd1 vssd1 vccd1 vccd1 _5824_/X sky130_fd_sc_hd__or3_1
XFILLER_22_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8543_ input3/X _8543_/D vssd1 vssd1 vccd1 vccd1 _8543_/Q sky130_fd_sc_hd__dfxtp_1
X_5755_ _5736_/A _5755_/B vssd1 vssd1 vccd1 vccd1 _5755_/X sky130_fd_sc_hd__and2b_1
X_8474_ input3/X _8474_/D vssd1 vssd1 vccd1 vccd1 _8474_/Q sky130_fd_sc_hd__dfxtp_1
X_4706_ _4706_/A _4706_/B _4706_/C vssd1 vssd1 vccd1 vccd1 _4707_/B sky130_fd_sc_hd__and3_1
X_5686_ _5686_/A _5800_/B vssd1 vssd1 vccd1 vccd1 _5689_/A sky130_fd_sc_hd__nand2_2
X_4637_ _4638_/A _4950_/A vssd1 vssd1 vccd1 vccd1 _4639_/A sky130_fd_sc_hd__and2_1
X_7425_ _8405_/A _8423_/B vssd1 vssd1 vccd1 vccd1 _8415_/A sky130_fd_sc_hd__and2_1
X_8659__75 vssd1 vssd1 vccd1 vccd1 _8659__75/HI _8768_/A sky130_fd_sc_hd__conb_1
XFILLER_89_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7356_ _7356_/A _7356_/B _7356_/C _7356_/D vssd1 vssd1 vccd1 vccd1 _7366_/B sky130_fd_sc_hd__and4_1
XFILLER_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4568_ _4570_/B _4568_/B _4568_/C vssd1 vssd1 vccd1 vccd1 _4569_/A sky130_fd_sc_hd__and3b_1
XFILLER_89_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7287_ _6822_/A _6822_/B _7286_/X vssd1 vssd1 vccd1 vccd1 _7288_/B sky130_fd_sc_hd__a21oi_2
X_6307_ _8529_/Q _8530_/Q _8533_/Q _6319_/D vssd1 vssd1 vccd1 vccd1 _6307_/X sky130_fd_sc_hd__o211a_1
X_4499_ _4689_/A vssd1 vssd1 vccd1 vccd1 _4510_/A sky130_fd_sc_hd__buf_2
X_6238_ _6238_/A _6238_/B vssd1 vssd1 vccd1 vccd1 _6239_/C sky130_fd_sc_hd__xnor2_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6169_ _6169_/A _6169_/B vssd1 vssd1 vccd1 vccd1 _6236_/C sky130_fd_sc_hd__xnor2_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5540_ _5540_/A vssd1 vssd1 vccd1 vccd1 _5664_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_8_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5471_ _5846_/A _5466_/Y _5829_/C vssd1 vssd1 vccd1 vccd1 _5472_/B sky130_fd_sc_hd__a21bo_1
X_7210_ _7187_/A _7187_/B _7187_/C vssd1 vssd1 vccd1 vccd1 _7211_/C sky130_fd_sc_hd__a21oi_1
X_4422_ _4713_/A vssd1 vssd1 vccd1 vccd1 _4438_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_8190_ _8190_/A _8190_/B _8190_/C vssd1 vssd1 vccd1 vccd1 _8191_/B sky130_fd_sc_hd__nor3_1
X_7141_ _7165_/B _7165_/A vssd1 vssd1 vccd1 vccd1 _7141_/X sky130_fd_sc_hd__and2b_1
X_4353_ _4357_/A vssd1 vssd1 vccd1 vccd1 _4353_/Y sky130_fd_sc_hd__inv_2
X_4284_ _4296_/A vssd1 vssd1 vccd1 vccd1 _4289_/A sky130_fd_sc_hd__clkbuf_2
X_7072_ _7121_/A _7070_/Y _7071_/X vssd1 vssd1 vccd1 vccd1 _7228_/A sky130_fd_sc_hd__a21o_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6023_ _6125_/A _6125_/B vssd1 vssd1 vccd1 vccd1 _6040_/A sky130_fd_sc_hd__xnor2_1
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7974_ _7974_/A _7974_/B vssd1 vssd1 vccd1 vccd1 _7975_/B sky130_fd_sc_hd__nor2_1
X_6925_ _6924_/A _6924_/C _6924_/B vssd1 vssd1 vccd1 vccd1 _6996_/B sky130_fd_sc_hd__a21o_1
XFILLER_81_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6856_ _6632_/A _6810_/A _6755_/B vssd1 vssd1 vccd1 vccd1 _6857_/B sky130_fd_sc_hd__o21a_1
XFILLER_50_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6787_ _6688_/A _6819_/B _6657_/A vssd1 vssd1 vccd1 vccd1 _6787_/X sky130_fd_sc_hd__a21o_1
XFILLER_50_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5807_ _5880_/A _5806_/X vssd1 vssd1 vccd1 vccd1 _5809_/B sky130_fd_sc_hd__or2b_1
X_8526_ input3/X _8526_/D vssd1 vssd1 vccd1 vccd1 _8526_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5738_ _5738_/A _6026_/A vssd1 vssd1 vccd1 vccd1 _5739_/A sky130_fd_sc_hd__or2_1
XFILLER_89_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8457_ input3/X _8457_/D vssd1 vssd1 vccd1 vccd1 _8457_/Q sky130_fd_sc_hd__dfxtp_4
X_5669_ _5669_/A _5669_/B _5669_/C vssd1 vssd1 vccd1 vccd1 _5669_/X sky130_fd_sc_hd__and3_1
X_7408_ _8565_/Q _7408_/B vssd1 vssd1 vccd1 vccd1 _7408_/X sky130_fd_sc_hd__or2_1
X_8388_ _8387_/Y _8426_/A _6462_/A vssd1 vssd1 vccd1 vccd1 _8388_/Y sky130_fd_sc_hd__a21oi_1
X_7339_ _7341_/B _7338_/C _7338_/A vssd1 vssd1 vccd1 vccd1 _7339_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_1_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_41 _8716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_52 _8772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_30 _8711_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_63 _8777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_74 _8786_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_85 _7613_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4971_ _5104_/C _5088_/B vssd1 vssd1 vccd1 vccd1 _5112_/D sky130_fd_sc_hd__or2_1
XFILLER_51_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6710_ _7079_/A vssd1 vssd1 vccd1 vccd1 _6947_/A sky130_fd_sc_hd__inv_2
X_7690_ _7690_/A _7690_/B vssd1 vssd1 vccd1 vccd1 _7691_/B sky130_fd_sc_hd__and2_1
X_6641_ _6739_/A vssd1 vssd1 vccd1 vccd1 _6643_/D sky130_fd_sc_hd__buf_2
X_6572_ _6570_/B _6570_/C _6513_/X vssd1 vssd1 vccd1 vccd1 _6714_/C sky130_fd_sc_hd__a21oi_2
X_8311_ _8311_/A _8311_/B vssd1 vssd1 vccd1 vccd1 _8344_/A sky130_fd_sc_hd__xnor2_1
X_5523_ _5426_/A _5648_/A _5406_/B _5522_/X vssd1 vssd1 vccd1 vccd1 _5540_/A sky130_fd_sc_hd__o31a_1
X_8242_ _8312_/B _8242_/B vssd1 vssd1 vccd1 vccd1 _8245_/A sky130_fd_sc_hd__xnor2_1
X_5454_ _6188_/A _5466_/A vssd1 vssd1 vccd1 vccd1 _5472_/A sky130_fd_sc_hd__nor2_1
X_4405_ _7575_/B vssd1 vssd1 vccd1 vccd1 _5178_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_5385_ _5385_/A _5385_/B vssd1 vssd1 vccd1 vccd1 _5563_/A sky130_fd_sc_hd__nand2_2
X_8629__45 vssd1 vssd1 vccd1 vccd1 _8629__45/HI _8724_/A sky130_fd_sc_hd__conb_1
X_8173_ _8173_/A _8085_/Y vssd1 vssd1 vccd1 vccd1 _8174_/B sky130_fd_sc_hd__or2b_1
X_7124_ _7149_/A _7149_/B vssd1 vssd1 vccd1 vccd1 _7126_/D sky130_fd_sc_hd__or2b_1
X_4336_ _4339_/A vssd1 vssd1 vccd1 vccd1 _4336_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7055_ _7055_/A _7055_/B vssd1 vssd1 vccd1 vccd1 _7109_/B sky130_fd_sc_hd__and2_1
X_4267_ _4270_/A vssd1 vssd1 vccd1 vccd1 _4267_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6006_ _6006_/A _6006_/B vssd1 vssd1 vccd1 vccd1 _6007_/B sky130_fd_sc_hd__and2_1
XFILLER_39_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7957_ _7944_/Y _7945_/X _7956_/X vssd1 vssd1 vccd1 vccd1 _7959_/A sky130_fd_sc_hd__a21boi_1
XFILLER_15_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6908_ _6889_/B _6905_/Y _6904_/A _6904_/Y vssd1 vssd1 vccd1 vccd1 _6909_/C sky130_fd_sc_hd__a211oi_2
X_7888_ _7888_/A _7888_/B vssd1 vssd1 vccd1 vccd1 _7888_/X sky130_fd_sc_hd__or2_1
X_6839_ _6839_/A _6839_/B vssd1 vssd1 vccd1 vccd1 _6840_/B sky130_fd_sc_hd__and2_1
XFILLER_24_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8509_ input3/X _8509_/D vssd1 vssd1 vccd1 vccd1 _8509_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5170_ _4973_/A _4898_/A _5089_/A _4975_/C _5153_/X vssd1 vssd1 vccd1 vccd1 _5171_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_68_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7811_ _7930_/A _7811_/B vssd1 vssd1 vccd1 vccd1 _7932_/B sky130_fd_sc_hd__and2_1
X_4954_ _5080_/B _5072_/A vssd1 vssd1 vccd1 vccd1 _4995_/C sky130_fd_sc_hd__or2_1
XFILLER_51_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7742_ _7742_/A _7885_/B _7885_/C vssd1 vssd1 vccd1 vccd1 _7861_/A sky130_fd_sc_hd__or3_2
XFILLER_17_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4885_ _4885_/A _5030_/C vssd1 vssd1 vccd1 vccd1 _5012_/C sky130_fd_sc_hd__or2_1
XFILLER_20_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7673_ _7672_/B _7672_/C _7678_/A vssd1 vssd1 vccd1 vccd1 _7674_/C sky130_fd_sc_hd__a21oi_1
X_6624_ _6745_/B vssd1 vssd1 vccd1 vccd1 _6977_/A sky130_fd_sc_hd__clkbuf_2
X_6555_ _6914_/A _6914_/C _6554_/Y vssd1 vssd1 vccd1 vccd1 _6929_/A sky130_fd_sc_hd__o21a_2
X_5506_ _5764_/B vssd1 vssd1 vccd1 vccd1 _5825_/B sky130_fd_sc_hd__clkbuf_2
X_6486_ _6486_/A _6486_/B vssd1 vssd1 vccd1 vccd1 _6506_/A sky130_fd_sc_hd__xnor2_2
X_8225_ _8227_/A _8225_/B vssd1 vssd1 vccd1 vccd1 _8225_/Y sky130_fd_sc_hd__nand2_1
X_5437_ _5437_/A _5437_/B vssd1 vssd1 vccd1 vccd1 _5459_/A sky130_fd_sc_hd__nor2_2
XFILLER_87_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5368_ _5526_/A _5368_/B _5368_/C vssd1 vssd1 vccd1 vccd1 _5370_/B sky130_fd_sc_hd__or3_1
X_8156_ _8156_/A _8276_/C vssd1 vssd1 vccd1 vccd1 _8277_/B sky130_fd_sc_hd__xnor2_1
X_4319_ _4320_/A vssd1 vssd1 vccd1 vccd1 _4319_/Y sky130_fd_sc_hd__inv_2
X_7107_ _7155_/A _7107_/B vssd1 vssd1 vccd1 vccd1 _7156_/A sky130_fd_sc_hd__xor2_1
X_8087_ _8037_/A _8037_/B _8038_/A _8086_/X vssd1 vssd1 vccd1 vccd1 _8171_/A sky130_fd_sc_hd__a31o_1
X_5299_ _8521_/Q vssd1 vssd1 vccd1 vccd1 _6270_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_74_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7038_ _7038_/A _7038_/B _7180_/B vssd1 vssd1 vccd1 vccd1 _7101_/A sky130_fd_sc_hd__nor3_2
XFILLER_59_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4670_ _4670_/A _4670_/B vssd1 vssd1 vccd1 vccd1 _4780_/B sky130_fd_sc_hd__nand2_1
X_6340_ _6340_/A vssd1 vssd1 vccd1 vccd1 _8530_/D sky130_fd_sc_hd__clkbuf_1
X_6271_ _6271_/A _6271_/B vssd1 vssd1 vccd1 vccd1 _6272_/B sky130_fd_sc_hd__nand2_1
X_5222_ _8494_/Q vssd1 vssd1 vccd1 vccd1 _6396_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_8010_ _8010_/A _8010_/B vssd1 vssd1 vccd1 vccd1 _8011_/B sky130_fd_sc_hd__or2_1
X_5153_ _5153_/A _5153_/B vssd1 vssd1 vccd1 vccd1 _5153_/X sky130_fd_sc_hd__or2_1
X_5084_ _5084_/A _5084_/B vssd1 vssd1 vccd1 vccd1 _5084_/X sky130_fd_sc_hd__or2_1
XFILLER_84_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8774_ _8774_/A _4367_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[21] sky130_fd_sc_hd__ebufn_8
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5986_ _6126_/A _5986_/B vssd1 vssd1 vccd1 vccd1 _5987_/B sky130_fd_sc_hd__xnor2_1
XFILLER_24_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4937_ _5138_/A _4937_/B vssd1 vssd1 vccd1 vccd1 _4937_/X sky130_fd_sc_hd__or2_1
X_7725_ _7725_/A _7725_/B _7725_/C vssd1 vssd1 vccd1 vccd1 _7841_/A sky130_fd_sc_hd__or3_1
X_4868_ _5074_/A _4993_/B vssd1 vssd1 vccd1 vccd1 _4868_/X sky130_fd_sc_hd__or2_1
XFILLER_20_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7656_ _7656_/A _7656_/B vssd1 vssd1 vccd1 vccd1 _7664_/A sky130_fd_sc_hd__xnor2_1
X_6607_ _6607_/A vssd1 vssd1 vccd1 vccd1 _6842_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4799_ _5050_/C _4913_/A vssd1 vssd1 vccd1 vccd1 _5020_/B sky130_fd_sc_hd__or2_2
X_7587_ _7899_/A _7587_/B vssd1 vssd1 vccd1 vccd1 _7677_/B sky130_fd_sc_hd__xor2_1
X_6538_ _6538_/A _8473_/Q vssd1 vssd1 vccd1 vccd1 _6539_/B sky130_fd_sc_hd__nor2_1
XFILLER_4_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6469_ _7410_/B _6468_/C _6538_/A vssd1 vssd1 vccd1 vccd1 _6470_/C sky130_fd_sc_hd__o21ai_1
X_8208_ _8210_/A _8213_/C vssd1 vssd1 vccd1 vccd1 _8209_/B sky130_fd_sc_hd__xor2_1
X_8139_ _8140_/A _8140_/B vssd1 vssd1 vccd1 vccd1 _8141_/A sky130_fd_sc_hd__nand2_1
XFILLER_75_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5840_ _5943_/A _5840_/B vssd1 vssd1 vccd1 vccd1 _5841_/B sky130_fd_sc_hd__xor2_2
X_5771_ _5824_/B _5824_/C vssd1 vssd1 vccd1 vccd1 _5772_/B sky130_fd_sc_hd__nor2_1
X_4722_ _4762_/A _4725_/A _4718_/A vssd1 vssd1 vccd1 vccd1 _4796_/A sky130_fd_sc_hd__or3b_4
X_8490_ input3/X _8490_/D vssd1 vssd1 vccd1 vccd1 _8490_/Q sky130_fd_sc_hd__dfxtp_1
X_7510_ _7805_/A _7921_/A vssd1 vssd1 vccd1 vccd1 _7546_/A sky130_fd_sc_hd__nand2_2
X_7441_ _8576_/Q vssd1 vssd1 vccd1 vccd1 _7766_/A sky130_fd_sc_hd__clkbuf_2
X_4653_ _5180_/A _4656_/S vssd1 vssd1 vccd1 vccd1 _4653_/Y sky130_fd_sc_hd__nor2_1
X_4584_ _4584_/A vssd1 vssd1 vccd1 vccd1 _5135_/A sky130_fd_sc_hd__buf_2
X_7372_ _7372_/A _7372_/B _7372_/C vssd1 vssd1 vccd1 vccd1 _7372_/X sky130_fd_sc_hd__or3_1
X_6323_ _6328_/B _7417_/A vssd1 vssd1 vccd1 vccd1 _7462_/A sky130_fd_sc_hd__or2_1
X_6254_ _6253_/B _6254_/B vssd1 vssd1 vccd1 vccd1 _6255_/B sky130_fd_sc_hd__and2b_1
X_5205_ _8480_/Q _5205_/B vssd1 vssd1 vccd1 vccd1 _5205_/X sky130_fd_sc_hd__or2_1
XFILLER_69_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6185_ _6104_/Y _6184_/Y _5984_/B vssd1 vssd1 vccd1 vccd1 _6186_/B sky130_fd_sc_hd__a21o_1
X_5136_ _5136_/A _5136_/B _5136_/C vssd1 vssd1 vccd1 vccd1 _5136_/X sky130_fd_sc_hd__or3_1
X_5067_ _5067_/A _5067_/B _5067_/C vssd1 vssd1 vccd1 vccd1 _5067_/X sky130_fd_sc_hd__or3_1
XFILLER_84_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8757_ _8757_/A _4343_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[4] sky130_fd_sc_hd__ebufn_8
X_5969_ _5923_/A _5923_/B _5924_/B _5924_/A vssd1 vssd1 vccd1 vccd1 _5993_/A sky130_fd_sc_hd__o2bb2ai_4
X_7708_ _8205_/B _7708_/B vssd1 vssd1 vccd1 vccd1 _7709_/A sky130_fd_sc_hd__nor2_1
X_8688_ _8688_/A _4264_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[5] sky130_fd_sc_hd__ebufn_8
XFILLER_32_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7639_ _7639_/A _7547_/B vssd1 vssd1 vccd1 vccd1 _7639_/X sky130_fd_sc_hd__or2b_1
XFILLER_75_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7990_ _8047_/A _7990_/B vssd1 vssd1 vccd1 vccd1 _7991_/B sky130_fd_sc_hd__and2_1
XFILLER_26_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6941_ _6941_/A _7152_/A vssd1 vssd1 vccd1 vccd1 _7055_/A sky130_fd_sc_hd__or2_1
XFILLER_47_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6872_ _7319_/A _6872_/B vssd1 vssd1 vccd1 vccd1 _6873_/B sky130_fd_sc_hd__xor2_2
XFILLER_34_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5823_ _5823_/A _5823_/B vssd1 vssd1 vccd1 vccd1 _5823_/Y sky130_fd_sc_hd__nand2_1
X_8542_ input3/X _8542_/D vssd1 vssd1 vccd1 vccd1 _8542_/Q sky130_fd_sc_hd__dfxtp_1
X_5754_ _5754_/A _5754_/B vssd1 vssd1 vccd1 vccd1 _5754_/X sky130_fd_sc_hd__or2_1
X_4705_ _4705_/A _4762_/C vssd1 vssd1 vccd1 vccd1 _4706_/C sky130_fd_sc_hd__nor2_1
X_8473_ input3/X _8473_/D vssd1 vssd1 vccd1 vccd1 _8473_/Q sky130_fd_sc_hd__dfxtp_1
X_5685_ _5685_/A _5860_/B _5685_/C vssd1 vssd1 vccd1 vccd1 _5691_/B sky130_fd_sc_hd__and3_1
X_4636_ _4949_/A _4640_/A _4635_/Y _4602_/X vssd1 vssd1 vccd1 vccd1 _8458_/D sky130_fd_sc_hd__o211a_1
XFILLER_8_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7424_ _8412_/B vssd1 vssd1 vccd1 vccd1 _8423_/B sky130_fd_sc_hd__clkbuf_1
X_7355_ _7350_/Y _7372_/B _7354_/Y vssd1 vssd1 vccd1 vccd1 _7356_/D sky130_fd_sc_hd__a21o_1
X_6306_ _8531_/Q vssd1 vssd1 vccd1 vccd1 _6319_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4567_ _8448_/Q _8449_/Q _4561_/B _8450_/Q vssd1 vssd1 vccd1 vccd1 _4568_/C sky130_fd_sc_hd__a31o_1
X_7286_ _7286_/A _7286_/B vssd1 vssd1 vccd1 vccd1 _7286_/X sky130_fd_sc_hd__and2_1
X_4498_ _6328_/A vssd1 vssd1 vccd1 vccd1 _4689_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6237_ _6236_/A _6236_/B _6236_/C vssd1 vssd1 vccd1 vccd1 _6239_/B sky130_fd_sc_hd__a21o_1
XFILLER_76_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6168_ _6168_/A _6168_/B vssd1 vssd1 vccd1 vccd1 _6169_/B sky130_fd_sc_hd__xor2_2
X_5119_ _5059_/A _5117_/X _5118_/X _5160_/A _5050_/A vssd1 vssd1 vccd1 vccd1 _5119_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6099_ _6046_/A _6046_/B _6098_/X vssd1 vssd1 vccd1 vccd1 _6174_/A sky130_fd_sc_hd__a21boi_1
XFILLER_17_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5470_ _5828_/A _6137_/A vssd1 vssd1 vccd1 vccd1 _5829_/C sky130_fd_sc_hd__or2_2
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4421_ _7498_/B vssd1 vssd1 vccd1 vccd1 _4713_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_8_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7140_ _7133_/A _7133_/B _7139_/X vssd1 vssd1 vccd1 vccd1 _7165_/A sky130_fd_sc_hd__a21bo_1
X_4352_ _4358_/A vssd1 vssd1 vccd1 vccd1 _4357_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_86_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4283_ _4283_/A vssd1 vssd1 vccd1 vccd1 _4283_/Y sky130_fd_sc_hd__inv_2
X_7071_ _7069_/A _6672_/A _7069_/B _6506_/A vssd1 vssd1 vccd1 vccd1 _7071_/X sky130_fd_sc_hd__o22a_1
XTAP_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6022_ _6124_/A _6124_/B vssd1 vssd1 vccd1 vccd1 _6125_/B sky130_fd_sc_hd__xor2_1
XFILLER_79_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7973_ _7974_/A _7974_/B vssd1 vssd1 vccd1 vccd1 _8046_/A sky130_fd_sc_hd__and2_2
XFILLER_81_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6924_ _6924_/A _6924_/B _6924_/C vssd1 vssd1 vccd1 vccd1 _6996_/A sky130_fd_sc_hd__nand3_4
XFILLER_35_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6855_ _7293_/A _7039_/B vssd1 vssd1 vccd1 vccd1 _6857_/A sky130_fd_sc_hd__nor2_1
XFILLER_22_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6786_ _7323_/A _6786_/B vssd1 vssd1 vccd1 vccd1 _6819_/B sky130_fd_sc_hd__or2_2
X_5806_ _5805_/A _5976_/A _5805_/D _5805_/C vssd1 vssd1 vccd1 vccd1 _5806_/X sky130_fd_sc_hd__a31o_1
X_5737_ _5488_/Y _5948_/A _5619_/B _5619_/A vssd1 vssd1 vccd1 vccd1 _5785_/A sky130_fd_sc_hd__a22o_1
X_8525_ input3/X _8525_/D vssd1 vssd1 vccd1 vccd1 _8525_/Q sky130_fd_sc_hd__dfxtp_1
X_8456_ input3/X _8456_/D vssd1 vssd1 vccd1 vccd1 _8456_/Q sky130_fd_sc_hd__dfxtp_1
X_7407_ _7403_/A _7406_/A _7406_/Y _6462_/X vssd1 vssd1 vccd1 vccd1 _8566_/D sky130_fd_sc_hd__a211o_1
X_5668_ _6075_/A _5668_/B vssd1 vssd1 vccd1 vccd1 _5669_/C sky130_fd_sc_hd__nor2_1
X_4619_ _4619_/A _4619_/B vssd1 vssd1 vccd1 vccd1 _4620_/A sky130_fd_sc_hd__nor2_1
X_5599_ _5599_/A _5599_/B vssd1 vssd1 vccd1 vccd1 _5600_/B sky130_fd_sc_hd__nand2_1
X_8387_ _8581_/Q vssd1 vssd1 vccd1 vccd1 _8387_/Y sky130_fd_sc_hd__inv_2
X_7338_ _7338_/A _7341_/B _7338_/C vssd1 vssd1 vccd1 vccd1 _7338_/X sky130_fd_sc_hd__and3_1
XFILLER_89_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7269_ _7030_/X _7268_/B _7268_/C _7268_/A vssd1 vssd1 vccd1 vccd1 _7270_/B sky130_fd_sc_hd__a211o_1
XFILLER_89_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_31 _8711_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_42 _8717_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_20 _8706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_75 _8786_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_53 _8772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_64 _8778_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_86 _7498_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4970_ _4970_/A _5035_/D vssd1 vssd1 vccd1 vccd1 _5088_/B sky130_fd_sc_hd__or2_1
X_6640_ _6640_/A _6640_/B _6964_/B vssd1 vssd1 vccd1 vccd1 _6739_/A sky130_fd_sc_hd__or3_1
XFILLER_32_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6571_ _6714_/B vssd1 vssd1 vccd1 vccd1 _6939_/B sky130_fd_sc_hd__clkbuf_2
X_8310_ _8310_/A _8310_/B vssd1 vssd1 vccd1 vccd1 _8311_/B sky130_fd_sc_hd__xnor2_1
X_5522_ _5522_/A _5427_/B vssd1 vssd1 vccd1 vccd1 _5522_/X sky130_fd_sc_hd__or2b_1
X_8241_ _8241_/A _8241_/B vssd1 vssd1 vccd1 vccd1 _8242_/B sky130_fd_sc_hd__xnor2_1
X_5453_ _5637_/A vssd1 vssd1 vccd1 vccd1 _5466_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4404_ _5180_/A _4404_/B _4655_/A vssd1 vssd1 vccd1 vccd1 _4469_/A sky130_fd_sc_hd__or3b_1
X_5384_ _5373_/A _5404_/B _5380_/X _5378_/X vssd1 vssd1 vccd1 vccd1 _5385_/B sky130_fd_sc_hd__a211o_1
X_8172_ _8085_/Y _8173_/A vssd1 vssd1 vccd1 vccd1 _8291_/A sky130_fd_sc_hd__nand2b_1
X_7123_ _7123_/A _7228_/A vssd1 vssd1 vccd1 vccd1 _7149_/B sky130_fd_sc_hd__xor2_1
X_4335_ _4339_/A vssd1 vssd1 vccd1 vccd1 _4335_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4266_ _4270_/A vssd1 vssd1 vccd1 vccd1 _4266_/Y sky130_fd_sc_hd__inv_2
X_7054_ _7054_/A _7116_/A vssd1 vssd1 vccd1 vccd1 _7055_/B sky130_fd_sc_hd__nand2_1
X_6005_ _6006_/A _6006_/B vssd1 vssd1 vccd1 vccd1 _6134_/A sky130_fd_sc_hd__nor2_1
XFILLER_55_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7956_ _7956_/A _7956_/B vssd1 vssd1 vccd1 vccd1 _7956_/X sky130_fd_sc_hd__xor2_1
X_6907_ _6907_/A _6907_/B vssd1 vssd1 vccd1 vccd1 _6909_/B sky130_fd_sc_hd__xnor2_1
X_7887_ _7886_/B _7886_/C _7886_/A vssd1 vssd1 vccd1 vccd1 _7898_/B sky130_fd_sc_hd__a21o_1
XFILLER_23_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6838_ _6838_/A _6838_/B vssd1 vssd1 vccd1 vccd1 _7325_/B sky130_fd_sc_hd__xor2_2
XFILLER_23_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6769_ _6823_/B _6769_/B vssd1 vssd1 vccd1 vccd1 _6771_/B sky130_fd_sc_hd__or2_1
X_8508_ input3/X _8508_/D vssd1 vssd1 vccd1 vccd1 _8508_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8439_ input3/X _8439_/D vssd1 vssd1 vccd1 vccd1 _8439_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7810_ _8176_/A _7810_/B _7830_/B vssd1 vssd1 vccd1 vccd1 _7811_/B sky130_fd_sc_hd__or3_1
XFILLER_36_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8790_ _8790_/A _4386_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[37] sky130_fd_sc_hd__ebufn_8
X_4953_ _4953_/A _4953_/B vssd1 vssd1 vccd1 vccd1 _5072_/A sky130_fd_sc_hd__nor2_1
XFILLER_51_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7741_ _7741_/A vssd1 vssd1 vccd1 vccd1 _7885_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_36_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7672_ _7678_/A _7672_/B _7672_/C vssd1 vssd1 vccd1 vccd1 _7796_/A sky130_fd_sc_hd__and3_1
X_4884_ _5099_/A _5026_/A _4957_/C _5033_/C vssd1 vssd1 vccd1 vccd1 _4884_/X sky130_fd_sc_hd__or4_1
X_6623_ _6623_/A _6623_/B vssd1 vssd1 vccd1 vccd1 _6745_/B sky130_fd_sc_hd__xnor2_4
XFILLER_20_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6554_ _7043_/A _6972_/A _6607_/A vssd1 vssd1 vccd1 vccd1 _6554_/Y sky130_fd_sc_hd__a21oi_2
X_6485_ _6714_/A _7183_/A vssd1 vssd1 vccd1 vccd1 _6505_/A sky130_fd_sc_hd__or2_1
X_5505_ _5602_/A _5505_/B vssd1 vssd1 vccd1 vccd1 _5516_/A sky130_fd_sc_hd__xnor2_1
XFILLER_10_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8224_ _8224_/A vssd1 vssd1 vccd1 vccd1 _8224_/Y sky130_fd_sc_hd__inv_2
X_5436_ _7554_/B _8522_/Q vssd1 vssd1 vccd1 vccd1 _5437_/B sky130_fd_sc_hd__and2b_1
XFILLER_87_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5367_ _5362_/C _5366_/X _5367_/S vssd1 vssd1 vccd1 vccd1 _5368_/C sky130_fd_sc_hd__mux2_1
X_8155_ _8274_/S _8155_/B vssd1 vssd1 vccd1 vccd1 _8276_/C sky130_fd_sc_hd__xnor2_1
X_4318_ _4320_/A vssd1 vssd1 vccd1 vccd1 _4318_/Y sky130_fd_sc_hd__inv_2
X_7106_ _7106_/A _7106_/B vssd1 vssd1 vccd1 vccd1 _7107_/B sky130_fd_sc_hd__xnor2_1
XFILLER_59_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8086_ _8086_/A _8086_/B vssd1 vssd1 vccd1 vccd1 _8086_/X sky130_fd_sc_hd__and2_1
X_5298_ _8522_/Q vssd1 vssd1 vccd1 vccd1 _6274_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_87_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7037_ _7037_/A vssd1 vssd1 vccd1 vccd1 _7180_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_47_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7939_ _7939_/A _7939_/B vssd1 vssd1 vccd1 vccd1 _7939_/Y sky130_fd_sc_hd__nand2_1
XFILLER_42_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6270_ _6270_/A _8507_/Q vssd1 vssd1 vccd1 vccd1 _6271_/B sky130_fd_sc_hd__or2b_1
XFILLER_88_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5221_ _8489_/Q _8488_/Q _6399_/A _6396_/B _8491_/Q vssd1 vssd1 vccd1 vccd1 _5221_/X
+ sky130_fd_sc_hd__a311o_1
X_5152_ _4935_/A _5020_/B _5146_/X _5151_/X vssd1 vssd1 vccd1 vccd1 _5152_/X sky130_fd_sc_hd__o31a_1
XFILLER_69_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5083_ _4974_/A _5064_/X _5160_/A vssd1 vssd1 vccd1 vccd1 _5084_/B sky130_fd_sc_hd__o21a_1
XFILLER_84_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8773_ _8773_/A _4366_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[20] sky130_fd_sc_hd__ebufn_8
XFILLER_64_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5985_ _5861_/A _5804_/B _6002_/A _5975_/X vssd1 vssd1 vccd1 vccd1 _5986_/B sky130_fd_sc_hd__a31oi_1
X_7724_ _7731_/A _7583_/A _7725_/C _7885_/A vssd1 vssd1 vccd1 vccd1 _7726_/B sky130_fd_sc_hd__o22ai_1
X_4936_ _4945_/A _5162_/B vssd1 vssd1 vccd1 vccd1 _4937_/B sky130_fd_sc_hd__or2_1
X_4867_ _5104_/C vssd1 vssd1 vccd1 vccd1 _5074_/A sky130_fd_sc_hd__clkbuf_2
X_7655_ _7655_/A _7655_/B _7547_/Y vssd1 vssd1 vccd1 vccd1 _7656_/B sky130_fd_sc_hd__or3b_2
X_6606_ _6606_/A vssd1 vssd1 vccd1 vccd1 _7033_/A sky130_fd_sc_hd__clkbuf_2
X_7586_ _7969_/A _7581_/Y _7952_/A vssd1 vssd1 vccd1 vccd1 _7587_/B sky130_fd_sc_hd__a21bo_1
X_4798_ _4899_/B _4798_/B vssd1 vssd1 vccd1 vccd1 _4913_/A sky130_fd_sc_hd__nor2_1
X_6537_ _8556_/Q _7644_/B vssd1 vssd1 vccd1 vccd1 _6539_/A sky130_fd_sc_hd__nor2_2
XFILLER_20_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6468_ _6538_/A _7410_/B _6468_/C vssd1 vssd1 vccd1 vccd1 _6470_/B sky130_fd_sc_hd__or3_1
X_6399_ _6399_/A _6399_/B _6399_/C _6399_/D vssd1 vssd1 vccd1 vccd1 _6424_/B sky130_fd_sc_hd__or4_4
X_5419_ _8514_/Q _7539_/B vssd1 vssd1 vccd1 vccd1 _5419_/Y sky130_fd_sc_hd__nand2_1
X_8207_ _8207_/A _8207_/B vssd1 vssd1 vccd1 vccd1 _8213_/C sky130_fd_sc_hd__xor2_1
X_8138_ _8054_/A _8366_/B _8326_/B vssd1 vssd1 vccd1 vccd1 _8140_/B sky130_fd_sc_hd__a21oi_1
XFILLER_87_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8069_ _8069_/A _8273_/A vssd1 vssd1 vccd1 vccd1 _8155_/B sky130_fd_sc_hd__nor2_1
XFILLER_47_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5770_ _5776_/A _5776_/B _5823_/B vssd1 vssd1 vccd1 vccd1 _5824_/C sky130_fd_sc_hd__a21oi_1
X_4721_ _5011_/A _5019_/B vssd1 vssd1 vccd1 vccd1 _4976_/A sky130_fd_sc_hd__or2_1
X_4652_ _5180_/A _4656_/S vssd1 vssd1 vccd1 vccd1 _4652_/X sky130_fd_sc_hd__and2_1
X_7440_ _7518_/A _7481_/B vssd1 vssd1 vccd1 vccd1 _7477_/A sky130_fd_sc_hd__nand2_1
X_4583_ _4945_/A vssd1 vssd1 vccd1 vccd1 _4584_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7371_ _6472_/X _8559_/Q _7362_/X _7370_/X vssd1 vssd1 vccd1 vccd1 _8559_/D sky130_fd_sc_hd__o22a_1
X_6322_ _6322_/A _6322_/B _6322_/C vssd1 vssd1 vccd1 vccd1 _7417_/A sky130_fd_sc_hd__and3_2
X_6253_ _6254_/B _6253_/B vssd1 vssd1 vccd1 vccd1 _6259_/B sky130_fd_sc_hd__and2b_1
X_5204_ _8578_/Q _5202_/X _5203_/X _5200_/X vssd1 vssd1 vccd1 vccd1 _8479_/D sky130_fd_sc_hd__o211a_1
XFILLER_88_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6184_ _6184_/A _6184_/B vssd1 vssd1 vccd1 vccd1 _6184_/Y sky130_fd_sc_hd__nand2_1
XFILLER_96_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5135_ _5135_/A _5135_/B _5135_/C vssd1 vssd1 vccd1 vccd1 _5135_/X sky130_fd_sc_hd__or3_1
XFILLER_69_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5066_ _5059_/X _5057_/X _5058_/X _5132_/A _4624_/A vssd1 vssd1 vccd1 vccd1 _5067_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_57_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8756_ _8756_/A _4345_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[3] sky130_fd_sc_hd__ebufn_8
X_5968_ _5959_/A _5959_/B _5967_/Y vssd1 vssd1 vccd1 vccd1 _6095_/B sky130_fd_sc_hd__a21o_1
XFILLER_40_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4919_ _5104_/D vssd1 vssd1 vccd1 vccd1 _5064_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_52_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7707_ _8371_/A _7707_/B vssd1 vssd1 vccd1 vccd1 _7708_/B sky130_fd_sc_hd__nor2_1
X_8687_ _8687_/A _4263_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[4] sky130_fd_sc_hd__ebufn_8
X_5899_ _6118_/A _5899_/B vssd1 vssd1 vccd1 vccd1 _5971_/A sky130_fd_sc_hd__nand2_1
XFILLER_32_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7638_ _7638_/A _7638_/B vssd1 vssd1 vccd1 vccd1 _7671_/A sky130_fd_sc_hd__and2_1
X_7569_ _7569_/A _7569_/B vssd1 vssd1 vccd1 vccd1 _7888_/A sky130_fd_sc_hd__xnor2_4
XFILLER_4_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6940_ _6940_/A vssd1 vssd1 vccd1 vccd1 _7152_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_54_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6871_ _6871_/A _6871_/B vssd1 vssd1 vccd1 vccd1 _6872_/B sky130_fd_sc_hd__nand2_1
XFILLER_62_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5822_ _5782_/A _5782_/B _5821_/Y vssd1 vssd1 vccd1 vccd1 _5925_/A sky130_fd_sc_hd__o21ai_2
X_8541_ input3/X _8541_/D vssd1 vssd1 vccd1 vccd1 _8541_/Q sky130_fd_sc_hd__dfxtp_1
X_5753_ _5754_/A _5754_/B vssd1 vssd1 vccd1 vccd1 _5753_/Y sky130_fd_sc_hd__nand2_1
XFILLER_34_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4704_ _4704_/A vssd1 vssd1 vccd1 vccd1 _8472_/D sky130_fd_sc_hd__clkbuf_1
X_8472_ input3/X _8472_/D vssd1 vssd1 vccd1 vccd1 _8472_/Q sky130_fd_sc_hd__dfxtp_1
X_5684_ _5684_/A vssd1 vssd1 vccd1 vccd1 _5860_/B sky130_fd_sc_hd__clkbuf_2
X_4635_ _4640_/A _5109_/A vssd1 vssd1 vccd1 vccd1 _4635_/Y sky130_fd_sc_hd__nand2_1
X_7423_ _8568_/Q vssd1 vssd1 vccd1 vccd1 _8412_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_7354_ _7354_/A _7354_/B vssd1 vssd1 vccd1 vccd1 _7354_/Y sky130_fd_sc_hd__xnor2_1
X_4566_ _8450_/Q _8449_/Q _4566_/C vssd1 vssd1 vccd1 vccd1 _4570_/B sky130_fd_sc_hd__and3_1
X_6305_ _8533_/Q vssd1 vssd1 vccd1 vccd1 _6351_/A sky130_fd_sc_hd__clkbuf_1
X_4497_ input2/X vssd1 vssd1 vccd1 vccd1 _6328_/A sky130_fd_sc_hd__clkbuf_2
X_7285_ _6839_/A _6838_/A _7284_/Y vssd1 vssd1 vccd1 vccd1 _7288_/A sky130_fd_sc_hd__o21ai_1
X_6236_ _6236_/A _6236_/B _6236_/C vssd1 vssd1 vccd1 vccd1 _6239_/A sky130_fd_sc_hd__nand3_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6167_ _6167_/A _6173_/B vssd1 vssd1 vccd1 vccd1 _6168_/B sky130_fd_sc_hd__xnor2_2
X_5118_ _5118_/A _5118_/B vssd1 vssd1 vccd1 vccd1 _5118_/X sky130_fd_sc_hd__or2_1
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6098_ _6098_/A _6045_/B vssd1 vssd1 vccd1 vccd1 _6098_/X sky130_fd_sc_hd__or2b_1
X_5049_ _5049_/A vssd1 vssd1 vccd1 vccd1 _5160_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_72_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8739_ _8739_/A _4326_/Y vssd1 vssd1 vccd1 vccd1 io_out[24] sky130_fd_sc_hd__ebufn_8
XFILLER_4_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4420_ _8468_/Q vssd1 vssd1 vccd1 vccd1 _7498_/B sky130_fd_sc_hd__buf_2
X_4351_ _4351_/A vssd1 vssd1 vccd1 vccd1 _4351_/Y sky130_fd_sc_hd__inv_2
X_4282_ _4283_/A vssd1 vssd1 vccd1 vccd1 _4282_/Y sky130_fd_sc_hd__inv_2
X_7070_ _7070_/A _7070_/B vssd1 vssd1 vccd1 vccd1 _7070_/Y sky130_fd_sc_hd__nand2_1
XTAP_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8664__80 vssd1 vssd1 vccd1 vccd1 _8664__80/HI _8773_/A sky130_fd_sc_hd__conb_1
X_6021_ _6021_/A _6021_/B vssd1 vssd1 vccd1 vccd1 _6124_/B sky130_fd_sc_hd__xnor2_1
XFILLER_67_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7972_ _7898_/A _7898_/B _7901_/B _7902_/B _7902_/A vssd1 vssd1 vccd1 vccd1 _7974_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6923_ _6899_/A _6899_/C _6899_/B vssd1 vssd1 vccd1 vccd1 _6924_/C sky130_fd_sc_hd__a21o_1
XFILLER_50_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6854_ _6854_/A _6854_/B vssd1 vssd1 vccd1 vccd1 _6860_/A sky130_fd_sc_hd__xor2_2
X_6785_ _7122_/C vssd1 vssd1 vccd1 vccd1 _7202_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_50_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5805_ _5805_/A _5976_/A _5805_/C _5805_/D vssd1 vssd1 vccd1 vccd1 _5880_/A sky130_fd_sc_hd__and4_1
XFILLER_50_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5736_ _5736_/A _5755_/B vssd1 vssd1 vccd1 vccd1 _5743_/A sky130_fd_sc_hd__xnor2_1
X_8524_ input3/X _8524_/D vssd1 vssd1 vccd1 vccd1 _8524_/Q sky130_fd_sc_hd__dfxtp_1
X_8455_ input3/X _8455_/D vssd1 vssd1 vccd1 vccd1 _8455_/Q sky130_fd_sc_hd__dfxtp_2
X_5667_ _5667_/A _5667_/B vssd1 vssd1 vccd1 vccd1 _5668_/B sky130_fd_sc_hd__and2_1
X_4618_ _5050_/A vssd1 vssd1 vccd1 vccd1 _5179_/A sky130_fd_sc_hd__buf_2
X_7406_ _7406_/A _7406_/B vssd1 vssd1 vccd1 vccd1 _7406_/Y sky130_fd_sc_hd__nor2_1
X_8386_ _8373_/X _8385_/X _6472_/X _8580_/Q vssd1 vssd1 vccd1 vccd1 _8580_/D sky130_fd_sc_hd__o2bb2a_1
X_5598_ _5599_/A _5599_/B vssd1 vssd1 vccd1 vccd1 _6084_/A sky130_fd_sc_hd__or2_1
X_7337_ _7337_/A _7337_/B vssd1 vssd1 vccd1 vccd1 _7356_/B sky130_fd_sc_hd__xnor2_2
XFILLER_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4549_ _8442_/Q _8443_/Q _4543_/B _8444_/Q vssd1 vssd1 vccd1 vccd1 _4550_/C sky130_fd_sc_hd__a31o_1
X_7268_ _7268_/A _7268_/B _7268_/C vssd1 vssd1 vccd1 vccd1 _7270_/A sky130_fd_sc_hd__nand3_1
XFILLER_89_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6219_ _6112_/A _6112_/B _6111_/A vssd1 vssd1 vccd1 vccd1 _6220_/B sky130_fd_sc_hd__a21o_1
X_7199_ _7201_/B _7201_/A vssd1 vssd1 vccd1 vccd1 _7200_/C sky130_fd_sc_hd__or2b_1
XINSDIODE2_10 _7358_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_43 _8717_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_21 _8706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_32 _8712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_65 _8778_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_76 _8787_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_54 _8773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6570_ _6570_/A _6570_/B _6570_/C vssd1 vssd1 vccd1 vccd1 _6714_/B sky130_fd_sc_hd__and3_1
X_5521_ _5521_/A _5521_/B vssd1 vssd1 vccd1 vccd1 _5554_/A sky130_fd_sc_hd__and2_1
XFILLER_8_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8240_ _8240_/A _8240_/B vssd1 vssd1 vccd1 vccd1 _8241_/B sky130_fd_sc_hd__xor2_1
X_5452_ _5778_/A vssd1 vssd1 vccd1 vccd1 _5637_/A sky130_fd_sc_hd__clkbuf_1
X_4403_ _7613_/B vssd1 vssd1 vccd1 vccd1 _4655_/A sky130_fd_sc_hd__clkbuf_1
X_8171_ _8171_/A _8171_/B vssd1 vssd1 vccd1 vccd1 _8173_/A sky130_fd_sc_hd__xor2_1
X_5383_ _5524_/A _5524_/B vssd1 vssd1 vccd1 vccd1 _5686_/A sky130_fd_sc_hd__xor2_4
X_7122_ _7202_/A _7185_/B _7122_/C _7070_/B vssd1 vssd1 vccd1 vccd1 _7149_/A sky130_fd_sc_hd__or4b_1
X_4334_ _4358_/A vssd1 vssd1 vccd1 vccd1 _4339_/A sky130_fd_sc_hd__clkbuf_4
X_7053_ _7105_/A _7045_/B _7033_/B vssd1 vssd1 vccd1 vccd1 _7109_/A sky130_fd_sc_hd__a21o_1
XFILLER_5_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4265_ _4390_/A vssd1 vssd1 vccd1 vccd1 _4270_/A sky130_fd_sc_hd__buf_2
X_6004_ _6004_/A _6004_/B vssd1 vssd1 vccd1 vccd1 _6006_/B sky130_fd_sc_hd__xnor2_1
XFILLER_55_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7955_ _8140_/A _7966_/A _8277_/A vssd1 vssd1 vccd1 vccd1 _7956_/B sky130_fd_sc_hd__o21ba_1
XFILLER_42_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6906_ _6904_/A _6904_/Y _6889_/B _6905_/Y vssd1 vssd1 vccd1 vccd1 _6909_/A sky130_fd_sc_hd__o211a_1
X_7886_ _7886_/A _7886_/B _7886_/C vssd1 vssd1 vccd1 vccd1 _7898_/A sky130_fd_sc_hd__nand3_1
X_6837_ _6837_/A _6848_/A vssd1 vssd1 vccd1 vccd1 _6838_/B sky130_fd_sc_hd__nand2_1
XFILLER_24_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6768_ _7054_/A _6768_/B vssd1 vssd1 vccd1 vccd1 _6769_/B sky130_fd_sc_hd__nor2_1
XFILLER_10_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8507_ input3/X _8507_/D vssd1 vssd1 vccd1 vccd1 _8507_/Q sky130_fd_sc_hd__dfxtp_1
X_6699_ _6698_/A _6698_/C _6698_/B vssd1 vssd1 vccd1 vccd1 _6700_/C sky130_fd_sc_hd__a21o_1
X_5719_ _5719_/A vssd1 vssd1 vccd1 vccd1 _5745_/A sky130_fd_sc_hd__inv_2
XFILLER_40_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8438_ input3/X _8438_/D vssd1 vssd1 vccd1 vccd1 _8438_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8369_ _8385_/A _8385_/B _8385_/C _8375_/B vssd1 vssd1 vccd1 vccd1 _8369_/X sky130_fd_sc_hd__or4_1
XFILLER_49_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8634__50 vssd1 vssd1 vccd1 vccd1 _8634__50/HI _8743_/A sky130_fd_sc_hd__conb_1
XFILLER_37_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4952_ _4893_/X _4932_/X _4949_/Y _5176_/S vssd1 vssd1 vccd1 vccd1 _4952_/X sky130_fd_sc_hd__a31o_1
X_7740_ _7740_/A vssd1 vssd1 vccd1 vccd1 _7885_/B sky130_fd_sc_hd__clkbuf_2
X_4883_ _5107_/C _4883_/B vssd1 vssd1 vccd1 vccd1 _5033_/C sky130_fd_sc_hd__or2_2
X_7671_ _7671_/A _7671_/B vssd1 vssd1 vccd1 vccd1 _7672_/C sky130_fd_sc_hd__or2_1
X_6622_ _6640_/A _6622_/B vssd1 vssd1 vccd1 vccd1 _6914_/B sky130_fd_sc_hd__nor2_1
XFILLER_32_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6553_ _6609_/A _6609_/B _6609_/C _6539_/A vssd1 vssd1 vccd1 vccd1 _6607_/A sky130_fd_sc_hd__a31o_1
X_6484_ _6939_/A vssd1 vssd1 vccd1 vccd1 _7183_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5504_ _5504_/A _5504_/B vssd1 vssd1 vccd1 vccd1 _5505_/B sky130_fd_sc_hd__xor2_1
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8223_ _8129_/A _8129_/B _8132_/A vssd1 vssd1 vccd1 vccd1 _8312_/B sky130_fd_sc_hd__o21ai_1
X_5435_ _8522_/Q _7554_/B vssd1 vssd1 vccd1 vccd1 _5437_/A sky130_fd_sc_hd__and2b_1
X_5366_ _5366_/A _5366_/B vssd1 vssd1 vccd1 vccd1 _5366_/X sky130_fd_sc_hd__or2_1
X_8154_ _8154_/A vssd1 vssd1 vccd1 vccd1 _8274_/S sky130_fd_sc_hd__clkbuf_2
X_4317_ _4320_/A vssd1 vssd1 vccd1 vccd1 _4317_/Y sky130_fd_sc_hd__inv_2
X_7105_ _7105_/A _7129_/A _7105_/C vssd1 vssd1 vccd1 vccd1 _7155_/A sky130_fd_sc_hd__nand3_2
XFILLER_59_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8085_ _8082_/A _8082_/B _8084_/Y vssd1 vssd1 vccd1 vccd1 _8085_/Y sky130_fd_sc_hd__a21oi_1
X_5297_ _8524_/Q vssd1 vssd1 vccd1 vccd1 _6286_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_7036_ _7044_/A _7044_/B _6745_/B vssd1 vssd1 vccd1 vccd1 _7036_/X sky130_fd_sc_hd__a21o_1
XFILLER_59_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7938_ _8184_/A _8184_/B _7937_/X vssd1 vssd1 vccd1 vccd1 _8016_/A sky130_fd_sc_hd__a21o_1
XFILLER_42_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7869_ _7869_/A _7869_/B vssd1 vssd1 vccd1 vccd1 _7870_/B sky130_fd_sc_hd__xnor2_2
XFILLER_50_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5220_ _8490_/Q vssd1 vssd1 vccd1 vccd1 _6396_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_5151_ _5151_/A _5151_/B _5151_/C _5151_/D vssd1 vssd1 vccd1 vccd1 _5151_/X sky130_fd_sc_hd__or4_1
XFILLER_69_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5082_ _5051_/A _5056_/C _5069_/X _5081_/X _5176_/S vssd1 vssd1 vccd1 vccd1 _5082_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_56_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8772_ _8772_/A _4365_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[19] sky130_fd_sc_hd__ebufn_8
XFILLER_64_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5984_ _5984_/A _5984_/B vssd1 vssd1 vccd1 vccd1 _6002_/A sky130_fd_sc_hd__nor2_2
X_7723_ _7888_/A _7740_/A _7741_/A vssd1 vssd1 vccd1 vccd1 _7747_/A sky130_fd_sc_hd__or3_2
XFILLER_40_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4935_ _4935_/A _4943_/B _5151_/B _5146_/A vssd1 vssd1 vccd1 vccd1 _4935_/X sky130_fd_sc_hd__or4_1
XFILLER_40_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4866_ _4866_/A vssd1 vssd1 vccd1 vccd1 _5104_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_32_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7654_ _7804_/A _7654_/B vssd1 vssd1 vccd1 vccd1 _7655_/B sky130_fd_sc_hd__nor2_1
X_4797_ _4880_/A _4881_/A vssd1 vssd1 vccd1 vccd1 _5050_/C sky130_fd_sc_hd__or2_2
X_6605_ _6623_/A _6623_/B vssd1 vssd1 vccd1 vccd1 _6606_/A sky130_fd_sc_hd__xor2_1
X_7585_ _7951_/A _8260_/A vssd1 vssd1 vccd1 vccd1 _7952_/A sky130_fd_sc_hd__or2_1
X_6536_ _6751_/B vssd1 vssd1 vccd1 vccd1 _6972_/A sky130_fd_sc_hd__buf_2
XFILLER_4_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6467_ _6455_/A _6452_/C _6459_/D _6466_/X vssd1 vssd1 vccd1 vccd1 _6468_/C sky130_fd_sc_hd__o31a_1
X_6398_ _6398_/A _6398_/B _6398_/C vssd1 vssd1 vccd1 vccd1 _6399_/D sky130_fd_sc_hd__or3_1
X_8206_ _8213_/D _8206_/B vssd1 vssd1 vccd1 vccd1 _8209_/A sky130_fd_sc_hd__nand2_1
X_5418_ _8514_/Q _7538_/B vssd1 vssd1 vccd1 vccd1 _5420_/A sky130_fd_sc_hd__nor2_1
X_5349_ _5349_/A _5349_/B vssd1 vssd1 vccd1 vccd1 _5349_/Y sky130_fd_sc_hd__nor2_1
X_8137_ _8066_/A _8135_/X _8136_/X vssd1 vssd1 vccd1 vccd1 _8247_/A sky130_fd_sc_hd__a21oi_1
XFILLER_87_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8068_ _7962_/A _7620_/A _8147_/B vssd1 vssd1 vccd1 vccd1 _8273_/A sky130_fd_sc_hd__a21o_1
X_7019_ _7019_/A _7019_/B _7019_/C _7019_/D vssd1 vssd1 vccd1 vccd1 _7019_/Y sky130_fd_sc_hd__nand4_4
XFILLER_47_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8604__20 vssd1 vssd1 vccd1 vccd1 _8604__20/HI _8699_/A sky130_fd_sc_hd__conb_1
XFILLER_59_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4720_ _4780_/A _4780_/B _4773_/A vssd1 vssd1 vccd1 vccd1 _5019_/B sky130_fd_sc_hd__nor3_2
X_4651_ _4651_/A vssd1 vssd1 vccd1 vccd1 _8461_/D sky130_fd_sc_hd__clkbuf_1
X_7370_ _7368_/Y _7369_/X _7366_/B vssd1 vssd1 vccd1 vccd1 _7370_/X sky130_fd_sc_hd__o21a_1
X_4582_ _8410_/A _4582_/B vssd1 vssd1 vccd1 vccd1 _8453_/D sky130_fd_sc_hd__nor2_1
X_6321_ _8546_/Q _6321_/B _8547_/Q _8545_/Q vssd1 vssd1 vccd1 vccd1 _6322_/C sky130_fd_sc_hd__and4b_1
X_6252_ _6246_/X _6251_/X _4668_/X _8516_/Q vssd1 vssd1 vccd1 vccd1 _8516_/D sky130_fd_sc_hd__o2bb2a_1
X_5203_ _8479_/Q _5205_/B vssd1 vssd1 vccd1 vccd1 _5203_/X sky130_fd_sc_hd__or2_1
XFILLER_88_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6183_ _6184_/A _6002_/A _6183_/S vssd1 vssd1 vccd1 vccd1 _6186_/A sky130_fd_sc_hd__mux2_1
X_5134_ _5020_/B _4842_/X _5059_/X _5132_/X _5133_/X vssd1 vssd1 vccd1 vccd1 _5134_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_69_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5065_ _5054_/X _5084_/A _5064_/X _4962_/X _5080_/A vssd1 vssd1 vccd1 vccd1 _5067_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_84_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8755_ _8755_/A _4348_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[2] sky130_fd_sc_hd__ebufn_8
XFILLER_12_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5967_ _5967_/A _5967_/B vssd1 vssd1 vccd1 vccd1 _5967_/Y sky130_fd_sc_hd__nor2_1
XFILLER_40_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4918_ _5020_/C _5074_/B vssd1 vssd1 vccd1 vccd1 _5104_/D sky130_fd_sc_hd__or2_1
X_8686_ _8686_/A _4262_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[3] sky130_fd_sc_hd__ebufn_8
XFILLER_52_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7706_ _7706_/A vssd1 vssd1 vccd1 vccd1 _8205_/B sky130_fd_sc_hd__inv_2
X_5898_ _5868_/A _5868_/B _5871_/A vssd1 vssd1 vccd1 vccd1 _5965_/A sky130_fd_sc_hd__a21bo_1
XFILLER_32_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7637_ _7637_/A _7637_/B vssd1 vssd1 vccd1 vccd1 _7638_/B sky130_fd_sc_hd__nand2_1
X_4849_ _5050_/C _4839_/X _4842_/X _4848_/X vssd1 vssd1 vccd1 vccd1 _4849_/X sky130_fd_sc_hd__o31a_1
XFILLER_20_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7568_ _7743_/A vssd1 vssd1 vccd1 vccd1 _7899_/A sky130_fd_sc_hd__clkbuf_2
X_6519_ _8564_/Q _8460_/Q vssd1 vssd1 vccd1 vccd1 _6563_/B sky130_fd_sc_hd__and2b_1
X_7499_ _7537_/A _7524_/B _7498_/X vssd1 vssd1 vccd1 vccd1 _7641_/A sky130_fd_sc_hd__a21o_2
XFILLER_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6870_ _6870_/A _6871_/A _6870_/C _6870_/D vssd1 vssd1 vccd1 vccd1 _6871_/B sky130_fd_sc_hd__nand4_1
XFILLER_22_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5821_ _5821_/A _5821_/B vssd1 vssd1 vccd1 vccd1 _5821_/Y sky130_fd_sc_hd__nand2_1
XFILLER_34_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8540_ input3/X _8540_/D vssd1 vssd1 vccd1 vccd1 _8540_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5752_ _5745_/A _5745_/B _5751_/X vssd1 vssd1 vccd1 vccd1 _5818_/A sky130_fd_sc_hd__a21o_1
X_4703_ _5370_/A _4703_/B _4703_/C vssd1 vssd1 vccd1 vccd1 _4704_/A sky130_fd_sc_hd__and3_1
X_8471_ input3/X _8471_/D vssd1 vssd1 vccd1 vccd1 _8471_/Q sky130_fd_sc_hd__dfxtp_1
X_5683_ _5683_/A _5683_/B vssd1 vssd1 vccd1 vccd1 _5811_/A sky130_fd_sc_hd__and2_1
X_4634_ _5125_/A vssd1 vssd1 vccd1 vccd1 _5109_/A sky130_fd_sc_hd__clkbuf_2
X_7422_ _7553_/A vssd1 vssd1 vccd1 vccd1 _8405_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7353_ _7359_/A _7352_/X _7254_/B vssd1 vssd1 vccd1 vccd1 _7372_/B sky130_fd_sc_hd__a21o_1
X_4565_ _8449_/Q _4566_/C _4564_/Y vssd1 vssd1 vccd1 vccd1 _8449_/D sky130_fd_sc_hd__a21oi_1
X_6304_ _8537_/Q vssd1 vssd1 vccd1 vccd1 _6362_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_4496_ _4496_/A vssd1 vssd1 vccd1 vccd1 _8735_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7284_ _6874_/A _6831_/B _6839_/A vssd1 vssd1 vccd1 vccd1 _7284_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_1_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6235_ _6235_/A _6235_/B vssd1 vssd1 vccd1 vccd1 _6235_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_69_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6166_ _6174_/A _6174_/B vssd1 vssd1 vccd1 vccd1 _6173_/B sky130_fd_sc_hd__xor2_1
X_5117_ _5117_/A _5117_/B _5117_/C vssd1 vssd1 vccd1 vccd1 _5117_/X sky130_fd_sc_hd__or3_1
XFILLER_84_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6097_ _5911_/A _5911_/B _5994_/B _5993_/B _5993_/A vssd1 vssd1 vccd1 vccd1 _6167_/A
+ sky130_fd_sc_hd__a32oi_4
X_5048_ _5046_/A _4864_/X _4952_/X _5047_/X vssd1 vssd1 vccd1 vccd1 _5048_/X sky130_fd_sc_hd__a31o_1
XFILLER_27_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8595__11 vssd1 vssd1 vccd1 vccd1 _8595__11/HI _8690_/A sky130_fd_sc_hd__conb_1
XFILLER_25_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8738_ _8738_/A _4325_/Y vssd1 vssd1 vccd1 vccd1 io_out[23] sky130_fd_sc_hd__ebufn_8
X_6999_ _6999_/A _6999_/B vssd1 vssd1 vccd1 vccd1 _7002_/A sky130_fd_sc_hd__xor2_2
XFILLER_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4350_ _4351_/A vssd1 vssd1 vccd1 vccd1 _4350_/Y sky130_fd_sc_hd__inv_2
X_4281_ _4283_/A vssd1 vssd1 vccd1 vccd1 _4281_/Y sky130_fd_sc_hd__inv_2
XTAP_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6020_ _6020_/A _6020_/B vssd1 vssd1 vccd1 vccd1 _6021_/B sky130_fd_sc_hd__nand2_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7971_ _8264_/A vssd1 vssd1 vccd1 vccd1 _7974_/A sky130_fd_sc_hd__inv_2
XFILLER_81_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6922_ _6983_/A _6983_/B vssd1 vssd1 vccd1 vccd1 _6924_/B sky130_fd_sc_hd__and2_1
X_6853_ _7297_/A _7297_/B vssd1 vssd1 vccd1 vccd1 _6854_/B sky130_fd_sc_hd__xor2_2
X_5804_ _5860_/B _5804_/B vssd1 vssd1 vccd1 vccd1 _5805_/D sky130_fd_sc_hd__or2_1
XFILLER_22_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6784_ _6784_/A vssd1 vssd1 vccd1 vccd1 _7122_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_22_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8523_ input3/X _8523_/D vssd1 vssd1 vccd1 vccd1 _8523_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5735_ _5735_/A _5735_/B vssd1 vssd1 vccd1 vccd1 _5755_/B sky130_fd_sc_hd__xnor2_1
X_8454_ input3/X _8454_/D vssd1 vssd1 vccd1 vccd1 _8454_/Q sky130_fd_sc_hd__dfxtp_1
X_5666_ _5667_/A _5667_/B vssd1 vssd1 vccd1 vccd1 _6075_/A sky130_fd_sc_hd__nor2_1
X_4617_ _4626_/B vssd1 vssd1 vccd1 vccd1 _5050_/A sky130_fd_sc_hd__clkbuf_2
X_7405_ _7405_/A _7405_/B vssd1 vssd1 vccd1 vccd1 _7406_/B sky130_fd_sc_hd__xnor2_1
X_8385_ _8385_/A _8385_/B _8385_/C _8385_/D vssd1 vssd1 vccd1 vccd1 _8385_/X sky130_fd_sc_hd__or4_1
X_5597_ _5594_/Y _5544_/B _5596_/X vssd1 vssd1 vccd1 vccd1 _5599_/B sky130_fd_sc_hd__a21oi_1
X_7336_ _7336_/A _7336_/B vssd1 vssd1 vccd1 vccd1 _7337_/B sky130_fd_sc_hd__xnor2_1
X_4548_ _8444_/Q _8443_/Q _4548_/C vssd1 vssd1 vccd1 vccd1 _4552_/B sky130_fd_sc_hd__and3_1
X_7267_ _7338_/A _7341_/B _7338_/C _7347_/A _7266_/Y vssd1 vssd1 vccd1 vccd1 _7268_/C
+ sky130_fd_sc_hd__a41o_1
XFILLER_89_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4479_ _4479_/A vssd1 vssd1 vccd1 vccd1 _8731_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_77_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6218_ _6134_/A _6133_/B _6131_/X vssd1 vssd1 vccd1 vccd1 _6220_/A sky130_fd_sc_hd__a21o_1
X_7198_ _7116_/A _7116_/B _7118_/B _7118_/A vssd1 vssd1 vccd1 vccd1 _7201_/A sky130_fd_sc_hd__a2bb2o_1
XINSDIODE2_33 _8712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_22 _8707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6149_ _5637_/B _5930_/B _6137_/C _6027_/B vssd1 vssd1 vccd1 vccd1 _6152_/A sky130_fd_sc_hd__a2bb2oi_1
XFILLER_38_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_11 _7372_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_77 _8787_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_55 _8773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_44 _8718_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_66 _8779_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5520_ _5520_/A _5520_/B vssd1 vssd1 vccd1 vccd1 _5521_/B sky130_fd_sc_hd__nand2_1
XFILLER_8_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5451_ _5774_/A vssd1 vssd1 vccd1 vccd1 _5778_/A sky130_fd_sc_hd__clkbuf_2
X_8170_ _8218_/B _8170_/B vssd1 vssd1 vccd1 vccd1 _8171_/B sky130_fd_sc_hd__xnor2_1
X_5382_ _5380_/X _5385_/A vssd1 vssd1 vccd1 vccd1 _5524_/B sky130_fd_sc_hd__and2b_2
X_4402_ _8463_/Q vssd1 vssd1 vccd1 vccd1 _7613_/B sky130_fd_sc_hd__buf_4
X_4333_ input1/X vssd1 vssd1 vccd1 vccd1 _4358_/A sky130_fd_sc_hd__clkbuf_2
X_7121_ _7121_/A _7121_/B vssd1 vssd1 vccd1 vccd1 _7185_/B sky130_fd_sc_hd__xnor2_2
X_7052_ _7052_/A _7052_/B vssd1 vssd1 vccd1 vccd1 _7114_/A sky130_fd_sc_hd__xnor2_1
XFILLER_59_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4264_ _4264_/A vssd1 vssd1 vccd1 vccd1 _4264_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6003_ _6104_/A _6177_/A vssd1 vssd1 vccd1 vccd1 _6004_/B sky130_fd_sc_hd__xor2_1
XFILLER_27_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7954_ _7954_/A _8260_/B vssd1 vssd1 vccd1 vccd1 _8277_/A sky130_fd_sc_hd__nor2_1
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6905_ _6888_/A _6888_/C _6888_/B vssd1 vssd1 vccd1 vccd1 _6905_/Y sky130_fd_sc_hd__o21ai_1
X_7885_ _7885_/A _7885_/B _7885_/C _8064_/A vssd1 vssd1 vccd1 vccd1 _7886_/C sky130_fd_sc_hd__or4_1
XFILLER_23_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6836_ _6836_/A _6837_/A _6836_/C vssd1 vssd1 vccd1 vccd1 _6848_/A sky130_fd_sc_hd__nand3_1
X_6767_ _6914_/A _6980_/B _6554_/Y vssd1 vssd1 vccd1 vccd1 _6768_/B sky130_fd_sc_hd__o21ai_1
X_8506_ input3/X _8506_/D vssd1 vssd1 vccd1 vccd1 _8506_/Q sky130_fd_sc_hd__dfxtp_1
X_5718_ _5718_/A _5718_/B vssd1 vssd1 vccd1 vccd1 _5749_/B sky130_fd_sc_hd__nand2_1
X_6698_ _6698_/A _6698_/B _6698_/C vssd1 vssd1 vccd1 vccd1 _6700_/B sky130_fd_sc_hd__nand3_1
X_5649_ _5649_/A _5795_/A vssd1 vssd1 vccd1 vccd1 _6053_/A sky130_fd_sc_hd__nor2_2
X_8437_ input3/X _8437_/D vssd1 vssd1 vccd1 vccd1 _8437_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8368_ _8370_/A _8366_/Y _8367_/X _7569_/B vssd1 vssd1 vccd1 vccd1 _8375_/B sky130_fd_sc_hd__o2bb2a_1
X_7319_ _7319_/A _6872_/B vssd1 vssd1 vccd1 vccd1 _7319_/X sky130_fd_sc_hd__or2b_1
XFILLER_77_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8299_ _8299_/A _8299_/B vssd1 vssd1 vccd1 vccd1 _8300_/B sky130_fd_sc_hd__xnor2_1
XFILLER_92_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4951_ _4951_/A vssd1 vssd1 vccd1 vccd1 _5176_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_64_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4882_ _4882_/A _5071_/A vssd1 vssd1 vccd1 vccd1 _4883_/B sky130_fd_sc_hd__and2_1
XFILLER_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7670_ _7671_/A _7671_/B vssd1 vssd1 vccd1 vccd1 _7672_/B sky130_fd_sc_hd__nand2_1
XFILLER_44_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6621_ _6733_/A _6620_/C _6829_/A vssd1 vssd1 vccd1 vccd1 _6645_/C sky130_fd_sc_hd__a21o_1
XFILLER_20_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6552_ _6972_/A _6913_/A vssd1 vssd1 vccd1 vccd1 _6914_/C sky130_fd_sc_hd__nor2_1
X_6483_ _7069_/A vssd1 vssd1 vccd1 vccd1 _6939_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_9_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5503_ _5625_/A _5625_/B vssd1 vssd1 vccd1 vccd1 _5504_/B sky130_fd_sc_hd__xor2_1
X_8222_ _8169_/A _8169_/B _8221_/X vssd1 vssd1 vccd1 vccd1 _8288_/A sky130_fd_sc_hd__a21o_1
X_5434_ _6281_/A _7553_/B vssd1 vssd1 vccd1 vccd1 _5461_/A sky130_fd_sc_hd__or2_1
X_8153_ _8276_/B vssd1 vssd1 vccd1 vccd1 _8156_/A sky130_fd_sc_hd__inv_2
X_7104_ _7103_/A _7103_/B _7103_/C vssd1 vssd1 vccd1 vccd1 _7105_/C sky130_fd_sc_hd__a21o_1
X_5365_ _8515_/Q vssd1 vssd1 vccd1 vccd1 _5526_/A sky130_fd_sc_hd__inv_2
X_4316_ _4320_/A vssd1 vssd1 vccd1 vccd1 _4316_/Y sky130_fd_sc_hd__inv_2
X_8084_ _8084_/A _8084_/B vssd1 vssd1 vccd1 vccd1 _8084_/Y sky130_fd_sc_hd__nor2_1
X_5296_ _8525_/Q vssd1 vssd1 vccd1 vccd1 _6293_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7035_ _7035_/A _7035_/B vssd1 vssd1 vccd1 vccd1 _7057_/A sky130_fd_sc_hd__xnor2_2
XFILLER_19_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7937_ _7936_/B _7937_/B vssd1 vssd1 vccd1 vccd1 _7937_/X sky130_fd_sc_hd__and2b_1
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7868_ _7868_/A _7875_/B vssd1 vssd1 vccd1 vccd1 _7869_/B sky130_fd_sc_hd__xnor2_1
X_6819_ _6819_/A _6819_/B vssd1 vssd1 vccd1 vccd1 _7286_/A sky130_fd_sc_hd__xor2_2
XFILLER_11_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7799_ _8205_/A _8371_/A _7707_/B _8213_/D vssd1 vssd1 vccd1 vccd1 _7800_/B sky130_fd_sc_hd__a31o_1
XFILLER_11_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5150_ _5132_/D _4937_/B _5147_/X _5148_/X _5156_/C vssd1 vssd1 vccd1 vccd1 _5151_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_69_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5081_ _5076_/X _5080_/X _4863_/X vssd1 vssd1 vccd1 vccd1 _5081_/X sky130_fd_sc_hd__a21o_1
XFILLER_37_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8771_ _8771_/A _4363_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[18] sky130_fd_sc_hd__ebufn_8
XFILLER_52_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5983_ _5983_/A _6101_/A vssd1 vssd1 vccd1 vccd1 _5987_/A sky130_fd_sc_hd__xnor2_1
X_4934_ _5147_/A vssd1 vssd1 vccd1 vccd1 _5146_/A sky130_fd_sc_hd__clkbuf_2
X_7722_ _7607_/B _7621_/A _7609_/B _7744_/A vssd1 vssd1 vccd1 vccd1 _7728_/A sky130_fd_sc_hd__a22o_1
X_4865_ _4968_/A vssd1 vssd1 vccd1 vccd1 _4987_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_32_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7653_ _7657_/A _7783_/B vssd1 vssd1 vccd1 vccd1 _7656_/A sky130_fd_sc_hd__xor2_1
X_4796_ _4796_/A _4796_/B vssd1 vssd1 vccd1 vccd1 _4881_/A sky130_fd_sc_hd__nor2_1
X_6604_ _6604_/A _6604_/B vssd1 vssd1 vccd1 vccd1 _6623_/B sky130_fd_sc_hd__and2_2
X_7584_ _7885_/A _7844_/A vssd1 vssd1 vccd1 vccd1 _8260_/A sky130_fd_sc_hd__xnor2_2
XFILLER_20_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6535_ _6751_/A vssd1 vssd1 vccd1 vccd1 _6914_/A sky130_fd_sc_hd__inv_2
X_6466_ _6466_/A _6466_/B vssd1 vssd1 vccd1 vccd1 _6466_/X sky130_fd_sc_hd__or2_1
X_8205_ _8205_/A _8205_/B _8206_/B vssd1 vssd1 vccd1 vccd1 _8361_/A sky130_fd_sc_hd__and3_1
X_6397_ _8499_/Q _8498_/Q _8506_/Q vssd1 vssd1 vccd1 vccd1 _6398_/C sky130_fd_sc_hd__or3_1
X_5417_ _5417_/A _5417_/B vssd1 vssd1 vccd1 vccd1 _6244_/A sky130_fd_sc_hd__nand2_2
X_5348_ _5341_/B _5343_/B _5341_/A vssd1 vssd1 vccd1 vccd1 _5349_/B sky130_fd_sc_hd__o21ba_1
X_8136_ _8136_/A _8136_/B vssd1 vssd1 vccd1 vccd1 _8136_/X sky130_fd_sc_hd__and2_1
X_8067_ _7956_/A _7956_/B _8277_/A vssd1 vssd1 vccd1 vccd1 _8073_/A sky130_fd_sc_hd__a21oi_1
X_7018_ _7017_/B _7017_/C _7017_/A vssd1 vssd1 vccd1 vccd1 _7019_/D sky130_fd_sc_hd__a21o_1
X_5279_ _5283_/C _5279_/B vssd1 vssd1 vccd1 vccd1 _8500_/D sky130_fd_sc_hd__nor2_1
XFILLER_75_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4650_ _4657_/B _4650_/B _4656_/S vssd1 vssd1 vccd1 vccd1 _4651_/A sky130_fd_sc_hd__and3_1
X_6320_ _6320_/A _6320_/B _6320_/C vssd1 vssd1 vccd1 vccd1 _6321_/B sky130_fd_sc_hd__and3_1
X_4581_ _8453_/Q _4575_/C _5322_/C vssd1 vssd1 vccd1 vccd1 _4582_/B sky130_fd_sc_hd__o21a_1
X_6251_ _6264_/B _6264_/C _6249_/Y _7399_/B vssd1 vssd1 vccd1 vccd1 _6251_/X sky130_fd_sc_hd__o31a_1
X_5202_ _5202_/A vssd1 vssd1 vccd1 vccd1 _5202_/X sky130_fd_sc_hd__clkbuf_2
X_6182_ _6182_/A _6182_/B vssd1 vssd1 vccd1 vccd1 _6215_/A sky130_fd_sc_hd__xnor2_1
X_5133_ _5179_/B _4900_/X _4904_/X _5092_/C vssd1 vssd1 vccd1 vccd1 _5133_/X sky130_fd_sc_hd__o22a_1
XFILLER_69_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5064_ _5064_/A _5064_/B _5064_/C _5064_/D vssd1 vssd1 vccd1 vccd1 _5064_/X sky130_fd_sc_hd__or4_1
XFILLER_72_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8754_ _8754_/A _4350_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[1] sky130_fd_sc_hd__ebufn_8
X_5966_ _5914_/A _5914_/B _5915_/A _5965_/X vssd1 vssd1 vccd1 vccd1 _6048_/A sky130_fd_sc_hd__a31o_1
X_4917_ _5099_/A vssd1 vssd1 vccd1 vccd1 _4955_/A sky130_fd_sc_hd__clkbuf_2
X_8685_ _8685_/A _4261_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[2] sky130_fd_sc_hd__ebufn_8
X_7705_ _8205_/A _7706_/A vssd1 vssd1 vccd1 vccd1 _8372_/A sky130_fd_sc_hd__xor2_1
XFILLER_12_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5897_ _5890_/A _5890_/B _5896_/X vssd1 vssd1 vccd1 vccd1 _5963_/A sky130_fd_sc_hd__a21oi_1
XFILLER_21_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4848_ _4848_/A _5132_/B _5132_/D _5051_/A vssd1 vssd1 vccd1 vccd1 _4848_/X sky130_fd_sc_hd__or4_1
X_7636_ _7637_/A _7637_/B vssd1 vssd1 vccd1 vccd1 _7638_/A sky130_fd_sc_hd__or2_1
XFILLER_20_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4779_ _4779_/A vssd1 vssd1 vccd1 vccd1 _4899_/A sky130_fd_sc_hd__clkbuf_2
X_7567_ _7594_/A _7594_/B _8367_/C vssd1 vssd1 vccd1 vccd1 _7743_/A sky130_fd_sc_hd__nand3_1
X_6518_ _7553_/B _8564_/Q vssd1 vssd1 vccd1 vccd1 _6575_/B sky130_fd_sc_hd__or2b_1
XFILLER_4_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7498_ _8571_/Q _7498_/B vssd1 vssd1 vccd1 vccd1 _7498_/X sky130_fd_sc_hd__and2b_1
X_6449_ _6445_/A _5294_/X _6432_/X _6448_/Y vssd1 vssd1 vccd1 vccd1 _8553_/D sky130_fd_sc_hd__a22o_1
X_8119_ _8120_/A _8120_/B vssd1 vssd1 vccd1 vccd1 _8233_/B sky130_fd_sc_hd__and2_1
XFILLER_87_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5820_ _5783_/A _5783_/B _5788_/A _5788_/B vssd1 vssd1 vccd1 vccd1 _5916_/A sky130_fd_sc_hd__a22oi_4
XFILLER_22_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5751_ _5744_/A _5751_/B vssd1 vssd1 vccd1 vccd1 _5751_/X sky130_fd_sc_hd__and2b_1
X_8470_ input3/X _8470_/D vssd1 vssd1 vccd1 vccd1 _8470_/Q sky130_fd_sc_hd__dfxtp_2
X_4702_ _7538_/B _4702_/B vssd1 vssd1 vccd1 vccd1 _4703_/C sky130_fd_sc_hd__or2_1
XFILLER_30_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5682_ _6249_/A _6259_/A _6249_/B vssd1 vssd1 vccd1 vccd1 _6264_/A sky130_fd_sc_hd__a21oi_1
X_7421_ _8584_/Q vssd1 vssd1 vccd1 vccd1 _7553_/A sky130_fd_sc_hd__inv_2
X_4633_ _4950_/A _4950_/B vssd1 vssd1 vccd1 vccd1 _5125_/A sky130_fd_sc_hd__or2_1
XFILLER_8_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7352_ _7352_/A _7352_/B vssd1 vssd1 vccd1 vccd1 _7352_/X sky130_fd_sc_hd__or2_1
X_4564_ _8449_/Q _4566_/C _4575_/A vssd1 vssd1 vccd1 vccd1 _4564_/Y sky130_fd_sc_hd__o21ai_1
X_6303_ _8542_/Q _8544_/Q _8543_/Q _8541_/Q vssd1 vssd1 vccd1 vccd1 _6320_/A sky130_fd_sc_hd__and4bb_1
X_7283_ _6862_/A _6862_/B _7282_/Y vssd1 vssd1 vccd1 vccd1 _7314_/A sky130_fd_sc_hd__a21oi_1
X_4495_ _8481_/Q _4495_/B vssd1 vssd1 vccd1 vccd1 _4496_/A sky130_fd_sc_hd__and2_1
X_6234_ _6238_/A _6238_/B _6090_/X vssd1 vssd1 vccd1 vccd1 _6235_/B sky130_fd_sc_hd__a21o_1
XFILLER_89_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6165_ _6224_/A _6165_/B vssd1 vssd1 vccd1 vccd1 _6174_/B sky130_fd_sc_hd__xor2_1
X_5116_ _5151_/A _5116_/B _5116_/C vssd1 vssd1 vccd1 vccd1 _5116_/X sky130_fd_sc_hd__or3_1
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6096_ _6048_/A _6048_/B _6095_/X vssd1 vssd1 vccd1 vccd1 _6168_/A sky130_fd_sc_hd__a21o_1
X_5047_ _4983_/X _5006_/X _5023_/X _5045_/X _5046_/Y vssd1 vssd1 vccd1 vccd1 _5047_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_27_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6998_ _6996_/X _6995_/Y _6994_/Y _6984_/X vssd1 vssd1 vccd1 vccd1 _7019_/B sky130_fd_sc_hd__o211ai_4
X_8737_ _8737_/A _4324_/Y vssd1 vssd1 vccd1 vccd1 io_out[22] sky130_fd_sc_hd__ebufn_8
XFILLER_13_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5949_ _5949_/A _6032_/B vssd1 vssd1 vccd1 vccd1 _5951_/A sky130_fd_sc_hd__xnor2_1
XFILLER_43_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7619_ _7618_/A _7618_/C _7618_/B vssd1 vssd1 vccd1 vccd1 _7741_/A sky130_fd_sc_hd__a21oi_1
XFILLER_21_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4280_ _4283_/A vssd1 vssd1 vccd1 vccd1 _4280_/Y sky130_fd_sc_hd__inv_2
XTAP_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7970_ _8142_/A _7888_/X _8319_/A vssd1 vssd1 vccd1 vccd1 _8264_/A sky130_fd_sc_hd__a21o_1
X_6921_ _6921_/A _6921_/B vssd1 vssd1 vccd1 vccd1 _6983_/B sky130_fd_sc_hd__xnor2_1
X_6852_ _6748_/B _6851_/Y _7291_/B vssd1 vssd1 vccd1 vccd1 _7297_/B sky130_fd_sc_hd__o21bai_2
X_5803_ _5918_/A _5803_/B vssd1 vssd1 vccd1 vccd1 _5805_/C sky130_fd_sc_hd__xnor2_1
XFILLER_22_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6783_ _6783_/A _6783_/B vssd1 vssd1 vccd1 vccd1 _7321_/A sky130_fd_sc_hd__xnor2_1
X_8522_ input3/X _8522_/D vssd1 vssd1 vccd1 vccd1 _8522_/Q sky130_fd_sc_hd__dfxtp_1
X_5734_ _5734_/A _5734_/B vssd1 vssd1 vccd1 vccd1 _5735_/B sky130_fd_sc_hd__xnor2_1
X_8453_ input3/X _8453_/D vssd1 vssd1 vccd1 vccd1 _8453_/Q sky130_fd_sc_hd__dfxtp_1
X_5665_ _5663_/Y _5664_/X _5539_/B _5548_/A vssd1 vssd1 vccd1 vccd1 _5667_/B sky130_fd_sc_hd__o31a_1
XFILLER_30_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4616_ _8456_/Q vssd1 vssd1 vccd1 vccd1 _4626_/B sky130_fd_sc_hd__inv_2
X_8384_ _8205_/A _8372_/A _8384_/S vssd1 vssd1 vccd1 vccd1 _8385_/D sky130_fd_sc_hd__mux2_1
X_7404_ _7404_/A _7408_/B vssd1 vssd1 vccd1 vccd1 _7405_/B sky130_fd_sc_hd__nand2_1
X_7335_ _7335_/A _7335_/B vssd1 vssd1 vccd1 vccd1 _7336_/B sky130_fd_sc_hd__xnor2_1
X_5596_ _6244_/A _5804_/B _5596_/C vssd1 vssd1 vccd1 vccd1 _5596_/X sky130_fd_sc_hd__and3_1
X_4547_ _8443_/Q _4548_/C _4546_/Y vssd1 vssd1 vccd1 vccd1 _8443_/D sky130_fd_sc_hd__a21oi_1
X_4478_ _8477_/Q _4480_/B vssd1 vssd1 vccd1 vccd1 _4479_/A sky130_fd_sc_hd__and2_1
X_7266_ _7171_/A _7265_/B _7263_/X vssd1 vssd1 vccd1 vccd1 _7266_/Y sky130_fd_sc_hd__a21oi_1
X_7197_ _7200_/B _7197_/B vssd1 vssd1 vccd1 vccd1 _7201_/B sky130_fd_sc_hd__nand2_1
X_6217_ _6122_/A _6122_/B _6216_/X vssd1 vssd1 vccd1 vccd1 _6221_/A sky130_fd_sc_hd__a21o_1
X_8655__71 vssd1 vssd1 vccd1 vccd1 _8655__71/HI _8764_/A sky130_fd_sc_hd__conb_1
XFILLER_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6148_ _6036_/A _6036_/B _6147_/X vssd1 vssd1 vccd1 vccd1 _6195_/A sky130_fd_sc_hd__a21bo_1
XINSDIODE2_23 _8707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_12 _7483_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_34 _8713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_45 _8718_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_67 _8779_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6079_ _6079_/A _6079_/B _6079_/C vssd1 vssd1 vccd1 vccd1 _6081_/A sky130_fd_sc_hd__nor3_1
XINSDIODE2_56 _8774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_78 _8788_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5450_ _8520_/Q _6482_/B vssd1 vssd1 vccd1 vccd1 _5774_/A sky130_fd_sc_hd__xnor2_4
X_4401_ _4949_/A _4593_/A _5180_/B vssd1 vssd1 vccd1 vccd1 _4404_/B sky130_fd_sc_hd__o21ai_1
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5381_ _8511_/Q _7501_/B vssd1 vssd1 vccd1 vccd1 _5385_/A sky130_fd_sc_hd__nand2_1
X_4332_ _4332_/A vssd1 vssd1 vccd1 vccd1 _4332_/Y sky130_fd_sc_hd__inv_2
X_7120_ _7070_/A _7070_/B _7071_/X vssd1 vssd1 vccd1 vccd1 _7121_/B sky130_fd_sc_hd__a21o_1
XFILLER_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7051_ _7052_/A _7052_/B vssd1 vssd1 vccd1 vccd1 _7064_/A sky130_fd_sc_hd__or2_1
X_4263_ _4264_/A vssd1 vssd1 vccd1 vccd1 _4263_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6002_ _6002_/A _6108_/B vssd1 vssd1 vccd1 vccd1 _6177_/A sky130_fd_sc_hd__xnor2_2
XFILLER_67_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7953_ _7886_/A _7886_/B _7886_/C vssd1 vssd1 vccd1 vccd1 _7966_/A sky130_fd_sc_hd__a21bo_1
XFILLER_39_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6904_ _6904_/A _6904_/B _6904_/C vssd1 vssd1 vccd1 vccd1 _6904_/Y sky130_fd_sc_hd__nor3_4
XFILLER_35_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7884_ _8317_/B _7885_/B _7885_/C _7950_/A _7961_/A vssd1 vssd1 vccd1 vccd1 _7886_/B
+ sky130_fd_sc_hd__o32ai_4
XFILLER_35_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6835_ _6858_/B _6834_/C _6929_/A vssd1 vssd1 vccd1 vccd1 _6836_/C sky130_fd_sc_hd__a21o_1
XFILLER_23_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6766_ _6914_/C vssd1 vssd1 vccd1 vccd1 _6980_/B sky130_fd_sc_hd__clkbuf_2
X_8505_ input3/X _8505_/D vssd1 vssd1 vccd1 vccd1 _8505_/Q sky130_fd_sc_hd__dfxtp_1
X_5717_ _5717_/A _5892_/B vssd1 vssd1 vccd1 vccd1 _6061_/A sky130_fd_sc_hd__xnor2_1
X_6697_ _7068_/B _6786_/B vssd1 vssd1 vccd1 vccd1 _6700_/A sky130_fd_sc_hd__nor2_1
X_8588__4 vssd1 vssd1 vccd1 vccd1 _8588__4/HI _8683_/A sky130_fd_sc_hd__conb_1
X_5648_ _5648_/A _5855_/B vssd1 vssd1 vccd1 vccd1 _5795_/A sky130_fd_sc_hd__or2_1
X_8436_ input3/X _8436_/D vssd1 vssd1 vccd1 vccd1 _8436_/Q sky130_fd_sc_hd__dfxtp_1
X_5579_ _5685_/A _5579_/B vssd1 vssd1 vccd1 vccd1 _5581_/A sky130_fd_sc_hd__nand2_1
X_8367_ _8367_/A _8367_/B _8367_/C vssd1 vssd1 vccd1 vccd1 _8367_/X sky130_fd_sc_hd__or3_1
X_7318_ _7318_/A _7318_/B vssd1 vssd1 vccd1 vccd1 _7332_/A sky130_fd_sc_hd__xor2_1
X_8298_ _8298_/A _8298_/B vssd1 vssd1 vccd1 vccd1 _8299_/B sky130_fd_sc_hd__nor2_1
X_7249_ _7351_/A _7351_/B vssd1 vssd1 vccd1 vccd1 _7352_/A sky130_fd_sc_hd__and2_1
XFILLER_49_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4950_ _4950_/A _4950_/B vssd1 vssd1 vccd1 vccd1 _4951_/A sky130_fd_sc_hd__nor2_1
X_4881_ _4881_/A vssd1 vssd1 vccd1 vccd1 _5071_/A sky130_fd_sc_hd__clkbuf_2
X_6620_ _6812_/A _6733_/A _6620_/C vssd1 vssd1 vccd1 vccd1 _6733_/B sky130_fd_sc_hd__nand3_1
XFILLER_20_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6551_ _6627_/A _6627_/B _6627_/C _6539_/A _6584_/A vssd1 vssd1 vccd1 vccd1 _6913_/A
+ sky130_fd_sc_hd__a311o_2
XFILLER_9_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5502_ _5502_/A _5624_/C vssd1 vssd1 vccd1 vccd1 _5625_/B sky130_fd_sc_hd__xnor2_1
X_6482_ _8561_/Q _6482_/B vssd1 vssd1 vccd1 vccd1 _7069_/A sky130_fd_sc_hd__xnor2_2
XFILLER_9_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5433_ _8460_/Q vssd1 vssd1 vccd1 vccd1 _7553_/B sky130_fd_sc_hd__clkbuf_4
X_8221_ _8168_/A _8221_/B vssd1 vssd1 vccd1 vccd1 _8221_/X sky130_fd_sc_hd__and2b_1
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8152_ _8152_/A _8152_/B vssd1 vssd1 vccd1 vccd1 _8159_/A sky130_fd_sc_hd__xor2_1
X_5364_ _5333_/X _5363_/Y _5360_/A _4511_/B vssd1 vssd1 vccd1 vccd1 _8514_/D sky130_fd_sc_hd__o2bb2a_1
X_4315_ _4327_/A vssd1 vssd1 vccd1 vccd1 _4320_/A sky130_fd_sc_hd__clkbuf_2
X_7103_ _7103_/A _7103_/B _7103_/C vssd1 vssd1 vccd1 vccd1 _7129_/A sky130_fd_sc_hd__nand3_2
X_5295_ _5293_/Y _5291_/C _5294_/X vssd1 vssd1 vccd1 vccd1 _8505_/D sky130_fd_sc_hd__a21boi_1
X_8083_ _8190_/A _8190_/B _8190_/C vssd1 vssd1 vccd1 vccd1 _8292_/A sky130_fd_sc_hd__o21a_1
X_7034_ _7033_/X _6975_/B _7034_/S vssd1 vssd1 vccd1 vccd1 _7035_/A sky130_fd_sc_hd__mux2_1
X_8625__41 vssd1 vssd1 vccd1 vccd1 _8625__41/HI _8720_/A sky130_fd_sc_hd__conb_1
XFILLER_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7936_ _7937_/B _7936_/B vssd1 vssd1 vccd1 vccd1 _8184_/B sky130_fd_sc_hd__xnor2_1
X_7867_ _7867_/A _7867_/B vssd1 vssd1 vccd1 vccd1 _7875_/B sky130_fd_sc_hd__xnor2_1
X_6818_ _7323_/A _7068_/B vssd1 vssd1 vccd1 vccd1 _6822_/A sky130_fd_sc_hd__nor2_1
XFILLER_23_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7798_ _7693_/A _7798_/B vssd1 vssd1 vccd1 vccd1 _8213_/D sky130_fd_sc_hd__and2b_1
X_6749_ _7043_/B _7038_/B _6748_/B vssd1 vssd1 vccd1 vccd1 _6749_/Y sky130_fd_sc_hd__o21bai_1
X_8419_ _8419_/A _8419_/B vssd1 vssd1 vccd1 vccd1 _8420_/A sky130_fd_sc_hd__and2_1
XFILLER_78_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5080_ _5080_/A _5080_/B _5080_/C _5080_/D vssd1 vssd1 vccd1 vccd1 _5080_/X sky130_fd_sc_hd__or4_1
XFILLER_56_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8770_ _8770_/A _4362_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[17] sky130_fd_sc_hd__ebufn_8
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5982_ _6104_/A _6102_/B vssd1 vssd1 vccd1 vccd1 _6101_/A sky130_fd_sc_hd__xor2_1
X_4933_ _4966_/A vssd1 vssd1 vccd1 vccd1 _5151_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_17_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7721_ _7623_/A _7623_/B _7720_/X vssd1 vssd1 vccd1 vccd1 _7738_/A sky130_fd_sc_hd__a21o_1
X_4864_ _4626_/A _4834_/X _4861_/X _5109_/A _4863_/X vssd1 vssd1 vccd1 vccd1 _4864_/X
+ sky130_fd_sc_hd__a2111o_1
X_7652_ _7658_/B _7652_/B vssd1 vssd1 vccd1 vccd1 _7783_/B sky130_fd_sc_hd__xnor2_2
X_4795_ _4875_/B _4796_/B vssd1 vssd1 vccd1 vccd1 _4880_/A sky130_fd_sc_hd__nor2_1
X_6603_ _6603_/A _7506_/B vssd1 vssd1 vccd1 vccd1 _6604_/B sky130_fd_sc_hd__nand2_1
X_7583_ _7583_/A vssd1 vssd1 vccd1 vccd1 _7844_/A sky130_fd_sc_hd__clkbuf_2
X_6534_ _6534_/A vssd1 vssd1 vccd1 vccd1 _6751_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_20_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6465_ _6465_/A vssd1 vssd1 vccd1 vccd1 _7410_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_5416_ _5900_/A _5408_/C _5685_/A vssd1 vssd1 vccd1 vccd1 _5429_/B sky130_fd_sc_hd__o21a_1
X_8204_ _8204_/A _8204_/B vssd1 vssd1 vccd1 vccd1 _8355_/A sky130_fd_sc_hd__nor2_1
X_6396_ _8491_/Q _6396_/B _8495_/Q _6396_/D vssd1 vssd1 vccd1 vccd1 _6398_/B sky130_fd_sc_hd__or4_1
X_5347_ _5347_/A _5347_/B vssd1 vssd1 vccd1 vccd1 _5349_/A sky130_fd_sc_hd__nor2_1
X_8135_ _8136_/A _8136_/B vssd1 vssd1 vccd1 vccd1 _8135_/X sky130_fd_sc_hd__or2_1
X_5278_ _8500_/Q _5276_/A _5264_/X vssd1 vssd1 vccd1 vccd1 _5279_/B sky130_fd_sc_hd__o21ai_1
X_8066_ _8066_/A _8066_/B vssd1 vssd1 vccd1 vccd1 _8074_/A sky130_fd_sc_hd__xnor2_1
X_7017_ _7017_/A _7017_/B _7017_/C vssd1 vssd1 vccd1 vccd1 _7019_/C sky130_fd_sc_hd__nand3_4
XFILLER_75_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7919_ _7984_/C vssd1 vssd1 vccd1 vccd1 _8249_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_62_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4580_ _5325_/B vssd1 vssd1 vccd1 vccd1 _5322_/C sky130_fd_sc_hd__clkbuf_2
X_6250_ _6328_/A vssd1 vssd1 vccd1 vccd1 _7399_/B sky130_fd_sc_hd__clkbuf_4
X_5201_ _8577_/Q _5188_/X _5199_/X _5200_/X vssd1 vssd1 vccd1 vccd1 _8478_/D sky130_fd_sc_hd__o211a_1
X_6181_ _6118_/A _6118_/B _6117_/B _6117_/A vssd1 vssd1 vccd1 vccd1 _6182_/B sky130_fd_sc_hd__o2bb2a_1
X_5132_ _5132_/A _5132_/B _5132_/C _5132_/D vssd1 vssd1 vccd1 vccd1 _5132_/X sky130_fd_sc_hd__or4_1
XFILLER_69_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5063_ _5087_/B _5080_/C _4848_/A vssd1 vssd1 vccd1 vccd1 _5084_/A sky130_fd_sc_hd__o21a_1
XFILLER_65_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8753_ _8753_/A _4387_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[0] sky130_fd_sc_hd__ebufn_8
X_5965_ _5965_/A _5965_/B vssd1 vssd1 vccd1 vccd1 _5965_/X sky130_fd_sc_hd__and2_1
X_4916_ _5104_/B _4989_/A _5030_/B vssd1 vssd1 vccd1 vccd1 _5164_/A sky130_fd_sc_hd__or3_1
XFILLER_80_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8684_ _8684_/A _4260_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[1] sky130_fd_sc_hd__ebufn_8
X_5896_ _5873_/A _5896_/B vssd1 vssd1 vccd1 vccd1 _5896_/X sky130_fd_sc_hd__and2b_1
X_7704_ _8371_/A _7707_/B vssd1 vssd1 vccd1 vccd1 _7706_/A sky130_fd_sc_hd__nand2_1
X_4847_ _4976_/A vssd1 vssd1 vccd1 vccd1 _5132_/D sky130_fd_sc_hd__clkbuf_2
X_7635_ _8317_/A _8052_/A _7635_/C _7969_/A vssd1 vssd1 vccd1 vccd1 _7637_/B sky130_fd_sc_hd__or4b_2
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4778_ _4960_/A vssd1 vssd1 vccd1 vccd1 _5132_/B sky130_fd_sc_hd__clkbuf_1
X_7566_ _7620_/A vssd1 vssd1 vccd1 vccd1 _8367_/C sky130_fd_sc_hd__inv_2
X_6517_ _6521_/A _6521_/B vssd1 vssd1 vccd1 vccd1 _6574_/B sky130_fd_sc_hd__or2_1
X_7497_ _8571_/Q _8468_/Q vssd1 vssd1 vccd1 vccd1 _7524_/B sky130_fd_sc_hd__xnor2_4
X_6448_ _6448_/A _6448_/B vssd1 vssd1 vccd1 vccd1 _6448_/Y sky130_fd_sc_hd__xnor2_1
X_6379_ _6380_/B _6380_/C _6378_/Y vssd1 vssd1 vccd1 vccd1 _8543_/D sky130_fd_sc_hd__a21oi_1
XFILLER_88_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8118_ _8105_/A _8305_/S _8123_/A _7925_/B vssd1 vssd1 vccd1 vccd1 _8120_/B sky130_fd_sc_hd__o22a_1
XFILLER_87_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8049_ _7976_/A _7976_/B _8048_/X vssd1 vssd1 vccd1 vccd1 _8077_/A sky130_fd_sc_hd__a21oi_1
XFILLER_56_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5750_ _6057_/A _6057_/B _5749_/X vssd1 vssd1 vccd1 vccd1 _5816_/B sky130_fd_sc_hd__a21o_1
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4701_ _7538_/B _4702_/B vssd1 vssd1 vccd1 vccd1 _4703_/B sky130_fd_sc_hd__nand2_1
X_5681_ _6083_/B _5681_/B vssd1 vssd1 vccd1 vccd1 _6249_/B sky130_fd_sc_hd__xnor2_1
X_4632_ _5441_/B _4862_/B vssd1 vssd1 vccd1 vccd1 _4950_/B sky130_fd_sc_hd__nor2_1
XFILLER_30_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7420_ _8397_/B _8391_/A _8584_/Q vssd1 vssd1 vccd1 vccd1 _7420_/X sky130_fd_sc_hd__o21a_1
X_7351_ _7351_/A _7351_/B vssd1 vssd1 vccd1 vccd1 _7352_/B sky130_fd_sc_hd__nor2_1
X_4563_ _4566_/C _4563_/B vssd1 vssd1 vccd1 vccd1 _8448_/D sky130_fd_sc_hd__nor2_1
X_4494_ _4494_/A vssd1 vssd1 vccd1 vccd1 _8734_/A sky130_fd_sc_hd__clkbuf_1
X_6302_ _8543_/Q vssd1 vssd1 vccd1 vccd1 _6380_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_7282_ _7282_/A _7282_/B vssd1 vssd1 vccd1 vccd1 _7282_/Y sky130_fd_sc_hd__nor2_1
XFILLER_89_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6233_ _6233_/A _6233_/B vssd1 vssd1 vccd1 vccd1 _6235_/A sky130_fd_sc_hd__xnor2_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6164_ _6223_/A _6164_/B vssd1 vssd1 vccd1 vccd1 _6165_/B sky130_fd_sc_hd__xnor2_1
X_5115_ _5099_/B _5058_/B _5088_/C _4584_/A vssd1 vssd1 vccd1 vccd1 _5116_/C sky130_fd_sc_hd__o31a_1
XFILLER_85_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6095_ _6047_/B _6095_/B vssd1 vssd1 vccd1 vccd1 _6095_/X sky130_fd_sc_hd__and2b_1
X_5046_ _5046_/A vssd1 vssd1 vccd1 vccd1 _5046_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6997_ _6984_/X _6994_/Y _6995_/Y _6996_/X vssd1 vssd1 vccd1 vccd1 _7019_/A sky130_fd_sc_hd__a211o_2
XFILLER_53_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8736_ _8736_/A _4323_/Y vssd1 vssd1 vccd1 vccd1 io_out[21] sky130_fd_sc_hd__ebufn_8
X_5948_ _5948_/A _6150_/A vssd1 vssd1 vccd1 vccd1 _6032_/B sky130_fd_sc_hd__nor2_1
XFILLER_40_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5879_ _6184_/A _5902_/A vssd1 vssd1 vccd1 vccd1 _5880_/C sky130_fd_sc_hd__nor2_1
X_7618_ _7618_/A _7618_/B _7618_/C vssd1 vssd1 vccd1 vccd1 _7740_/A sky130_fd_sc_hd__and3_1
XFILLER_5_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7549_ _7549_/A _7549_/B vssd1 vssd1 vccd1 vccd1 _7677_/A sky130_fd_sc_hd__xnor2_1
XFILLER_4_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6920_ _6977_/A _6978_/A _6977_/B vssd1 vssd1 vccd1 vccd1 _6921_/B sky130_fd_sc_hd__o21ba_1
XFILLER_54_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6851_ _7293_/A _6977_/B vssd1 vssd1 vccd1 vccd1 _6851_/Y sky130_fd_sc_hd__nor2_1
XFILLER_35_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5802_ _5689_/A _6126_/A _5801_/Y vssd1 vssd1 vccd1 vccd1 _5803_/B sky130_fd_sc_hd__o21a_1
XFILLER_35_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6782_ _7328_/A _7279_/A vssd1 vssd1 vccd1 vccd1 _6783_/B sky130_fd_sc_hd__nand2_1
XFILLER_50_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8521_ input3/X _8521_/D vssd1 vssd1 vccd1 vccd1 _8521_/Q sky130_fd_sc_hd__dfxtp_1
X_5733_ _5948_/A _5733_/B vssd1 vssd1 vccd1 vccd1 _5734_/B sky130_fd_sc_hd__nor2_1
X_5664_ _5664_/A _5664_/B vssd1 vssd1 vccd1 vccd1 _5664_/X sky130_fd_sc_hd__and2_1
XFILLER_30_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8452_ input3/X _8452_/D vssd1 vssd1 vccd1 vccd1 _8452_/Q sky130_fd_sc_hd__dfxtp_1
X_4615_ _5174_/S _4643_/A vssd1 vssd1 vccd1 vccd1 _4629_/A sky130_fd_sc_hd__nand2_1
X_7403_ _7403_/A _7403_/B vssd1 vssd1 vccd1 vccd1 _7408_/B sky130_fd_sc_hd__or2_1
X_8383_ _8373_/X _8382_/X _6261_/X _8579_/Q vssd1 vssd1 vccd1 vccd1 _8579_/D sky130_fd_sc_hd__o2bb2a_1
X_5595_ _5650_/A vssd1 vssd1 vccd1 vccd1 _5804_/B sky130_fd_sc_hd__clkbuf_2
X_7334_ _7334_/A _7334_/B vssd1 vssd1 vccd1 vccd1 _7335_/B sky130_fd_sc_hd__xnor2_1
X_4546_ _8443_/Q _4548_/C _4536_/X vssd1 vssd1 vccd1 vccd1 _4546_/Y sky130_fd_sc_hd__o21ai_1
X_7265_ _7263_/X _7265_/B vssd1 vssd1 vccd1 vccd1 _7347_/A sky130_fd_sc_hd__and2b_1
X_4477_ _4477_/A vssd1 vssd1 vccd1 vccd1 _8730_/A sky130_fd_sc_hd__clkbuf_1
X_7196_ _7196_/A _7196_/B _7196_/C vssd1 vssd1 vccd1 vccd1 _7197_/B sky130_fd_sc_hd__or3_1
X_6216_ _6119_/B _6216_/B vssd1 vssd1 vccd1 vccd1 _6216_/X sky130_fd_sc_hd__and2b_1
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6147_ _6147_/A _6154_/B vssd1 vssd1 vccd1 vccd1 _6147_/X sky130_fd_sc_hd__or2b_1
XFILLER_38_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_13 _7483_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_24 _8708_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_35 _8713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_57 _8774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6078_ _6078_/A _6078_/B _6078_/C vssd1 vssd1 vccd1 vccd1 _6079_/C sky130_fd_sc_hd__nor3_1
XINSDIODE2_68 _8780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8670__86 vssd1 vssd1 vccd1 vccd1 _8670__86/HI _8779_/A sky130_fd_sc_hd__conb_1
XINSDIODE2_46 _8743_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_79 _8788_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5029_ _5055_/A vssd1 vssd1 vccd1 vccd1 _5099_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_38_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8719_ _8719_/A _4301_/Y vssd1 vssd1 vccd1 vccd1 io_out[4] sky130_fd_sc_hd__ebufn_8
XFILLER_70_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4400_ _6521_/B vssd1 vssd1 vccd1 vccd1 _5180_/B sky130_fd_sc_hd__clkbuf_1
X_5380_ _8511_/Q _5380_/B vssd1 vssd1 vccd1 vccd1 _5380_/X sky130_fd_sc_hd__and2b_1
X_4331_ _4332_/A vssd1 vssd1 vccd1 vccd1 _4331_/Y sky130_fd_sc_hd__inv_2
X_7050_ _7050_/A _7050_/B vssd1 vssd1 vccd1 vccd1 _7052_/B sky130_fd_sc_hd__xnor2_2
X_4262_ _4264_/A vssd1 vssd1 vccd1 vccd1 _4262_/Y sky130_fd_sc_hd__inv_2
X_6001_ _5694_/A _5861_/C _6126_/B vssd1 vssd1 vccd1 vccd1 _6108_/B sky130_fd_sc_hd__mux2_1
XFILLER_79_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7952_ _7952_/A _8053_/B _7952_/C vssd1 vssd1 vccd1 vccd1 _8140_/A sky130_fd_sc_hd__and3_1
XFILLER_39_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6903_ _6883_/X _6900_/Y _6924_/A _6895_/Y vssd1 vssd1 vccd1 vccd1 _6904_/C sky130_fd_sc_hd__o211a_1
X_7883_ _7945_/A vssd1 vssd1 vccd1 vccd1 _8142_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_62_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6834_ _6929_/A _6858_/B _6834_/C vssd1 vssd1 vccd1 vccd1 _6837_/A sky130_fd_sc_hd__nand3_1
X_6765_ _7118_/A _6929_/A vssd1 vssd1 vccd1 vccd1 _6823_/B sky130_fd_sc_hd__nor2_1
XFILLER_50_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8504_ input3/X _8504_/D vssd1 vssd1 vccd1 vccd1 _8504_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5716_ _5889_/A _5716_/B vssd1 vssd1 vccd1 vccd1 _5892_/B sky130_fd_sc_hd__nand2_1
X_6696_ _6675_/A _6674_/C _6780_/A vssd1 vssd1 vccd1 vccd1 _6698_/C sky130_fd_sc_hd__a21o_1
XFILLER_40_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8435_ input3/X _8435_/D vssd1 vssd1 vccd1 vccd1 _8435_/Q sky130_fd_sc_hd__dfxtp_1
X_5647_ _5528_/B _5530_/B _5646_/Y vssd1 vssd1 vccd1 vccd1 _5855_/B sky130_fd_sc_hd__a21o_1
XFILLER_40_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8366_ _8366_/A _8366_/B vssd1 vssd1 vccd1 vccd1 _8366_/Y sky130_fd_sc_hd__nand2_1
X_5578_ _5578_/A _5578_/B vssd1 vssd1 vccd1 vccd1 _6248_/A sky130_fd_sc_hd__xnor2_2
X_7317_ _6569_/B _6819_/B _6569_/A vssd1 vssd1 vccd1 vccd1 _7318_/B sky130_fd_sc_hd__o21ba_1
X_8297_ _8287_/A _8297_/B vssd1 vssd1 vccd1 vccd1 _8298_/B sky130_fd_sc_hd__and2b_1
X_4529_ _4533_/C _4529_/B vssd1 vssd1 vccd1 vccd1 _8437_/D sky130_fd_sc_hd__nor2_1
X_7248_ _7248_/A _7248_/B _7250_/B vssd1 vssd1 vccd1 vccd1 _7351_/B sky130_fd_sc_hd__and3_1
XFILLER_49_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7179_ _7038_/A _7175_/B _6977_/B _7180_/A vssd1 vssd1 vccd1 vccd1 _7180_/C sky130_fd_sc_hd__o22a_1
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4880_ _4880_/A vssd1 vssd1 vccd1 vccd1 _5107_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_51_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6550_ _6609_/C vssd1 vssd1 vccd1 vccd1 _6627_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5501_ _5774_/A _5764_/B _5764_/C vssd1 vssd1 vccd1 vccd1 _5624_/C sky130_fd_sc_hd__or3_2
X_6481_ _6481_/A vssd1 vssd1 vccd1 vccd1 _6714_/A sky130_fd_sc_hd__clkbuf_2
X_8220_ _8034_/A _8034_/B _8115_/B _8114_/B _8114_/A vssd1 vssd1 vccd1 vccd1 _8346_/A
+ sky130_fd_sc_hd__a32oi_4
X_5432_ _5497_/A _5432_/B vssd1 vssd1 vccd1 vccd1 _5445_/A sky130_fd_sc_hd__and2_1
X_8151_ _7756_/B _8063_/B _8064_/B _8064_/A vssd1 vssd1 vccd1 vccd1 _8152_/B sky130_fd_sc_hd__o22a_1
X_5363_ _5363_/A _5363_/B vssd1 vssd1 vccd1 vccd1 _5363_/Y sky130_fd_sc_hd__nand2_1
X_4314_ _4314_/A vssd1 vssd1 vccd1 vccd1 _4314_/Y sky130_fd_sc_hd__inv_2
X_7102_ _7102_/A _7102_/B vssd1 vssd1 vccd1 vccd1 _7103_/C sky130_fd_sc_hd__xnor2_1
XFILLER_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5294_ _5294_/A vssd1 vssd1 vccd1 vccd1 _5294_/X sky130_fd_sc_hd__clkbuf_4
X_8082_ _8082_/A _8082_/B vssd1 vssd1 vccd1 vccd1 _8190_/C sky130_fd_sc_hd__xor2_1
X_7033_ _7033_/A _7033_/B _7044_/B vssd1 vssd1 vccd1 vccd1 _7033_/X sky130_fd_sc_hd__or3b_2
XFILLER_95_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8640__56 vssd1 vssd1 vccd1 vccd1 _8640__56/HI _8749_/A sky130_fd_sc_hd__conb_1
X_8590__6 vssd1 vssd1 vccd1 vccd1 _8590__6/HI _8685_/A sky130_fd_sc_hd__conb_1
XFILLER_82_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7935_ _7935_/A _7935_/B vssd1 vssd1 vccd1 vccd1 _7936_/B sky130_fd_sc_hd__xnor2_1
XFILLER_35_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7866_ _7866_/A _7866_/B vssd1 vssd1 vccd1 vccd1 _7867_/B sky130_fd_sc_hd__xnor2_2
XFILLER_35_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6817_ _6826_/A _6817_/B _6817_/C vssd1 vssd1 vccd1 vccd1 _6870_/A sky130_fd_sc_hd__nand3_1
XFILLER_51_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7797_ _8210_/A _8213_/B vssd1 vssd1 vccd1 vccd1 _8206_/B sky130_fd_sc_hd__nor2b_1
XFILLER_23_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6748_ _7038_/B _6748_/B vssd1 vssd1 vccd1 vccd1 _7291_/B sky130_fd_sc_hd__and2b_1
X_6679_ _6939_/A _6679_/B vssd1 vssd1 vccd1 vccd1 _6690_/C sky130_fd_sc_hd__nor2_1
X_8418_ _8417_/X _8428_/A _8418_/S vssd1 vssd1 vccd1 vccd1 _8419_/B sky130_fd_sc_hd__mux2_1
X_8349_ _8345_/X _8346_/X _8348_/X vssd1 vssd1 vccd1 vccd1 _8349_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_78_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5981_ _5984_/B _5981_/B _6106_/B vssd1 vssd1 vccd1 vccd1 _6102_/B sky130_fd_sc_hd__and3b_1
X_4932_ _5067_/A _4932_/B _4932_/C vssd1 vssd1 vccd1 vccd1 _4932_/X sky130_fd_sc_hd__or3_1
X_7720_ _7635_/C _7720_/B vssd1 vssd1 vccd1 vccd1 _7720_/X sky130_fd_sc_hd__and2b_1
X_7651_ _7769_/A _7660_/A vssd1 vssd1 vccd1 vccd1 _7652_/B sky130_fd_sc_hd__xnor2_1
X_4863_ _4863_/A vssd1 vssd1 vccd1 vccd1 _4863_/X sky130_fd_sc_hd__clkbuf_2
X_6602_ _6500_/A _6500_/B _6499_/A vssd1 vssd1 vccd1 vccd1 _6623_/A sky130_fd_sc_hd__a21oi_4
XFILLER_32_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4794_ _5055_/A _5018_/A vssd1 vssd1 vccd1 vccd1 _4914_/A sky130_fd_sc_hd__or2_1
X_7582_ _7607_/A vssd1 vssd1 vccd1 vccd1 _7885_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_32_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6533_ _7054_/A _6721_/A _6679_/B vssd1 vssd1 vccd1 vccd1 _7093_/A sky130_fd_sc_hd__o21a_2
X_6464_ _8556_/Q vssd1 vssd1 vccd1 vccd1 _6538_/A sky130_fd_sc_hd__inv_2
XFILLER_21_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5415_ _5579_/B vssd1 vssd1 vccd1 vccd1 _5900_/A sky130_fd_sc_hd__clkbuf_2
X_8203_ _8202_/A _8202_/C _8202_/B vssd1 vssd1 vccd1 vccd1 _8204_/B sky130_fd_sc_hd__o21a_1
X_6395_ _8489_/Q _8488_/Q vssd1 vssd1 vccd1 vccd1 _6398_/A sky130_fd_sc_hd__nand2_1
X_5346_ _8512_/Q _5360_/B vssd1 vssd1 vccd1 vccd1 _5347_/B sky130_fd_sc_hd__and2b_1
X_8134_ _8076_/A _8134_/B vssd1 vssd1 vccd1 vccd1 _8165_/B sky130_fd_sc_hd__and2b_1
X_5277_ _8500_/Q _8499_/Q _5277_/C vssd1 vssd1 vccd1 vccd1 _5283_/C sky130_fd_sc_hd__and3_1
X_8065_ _8136_/A _8136_/B vssd1 vssd1 vccd1 vccd1 _8066_/B sky130_fd_sc_hd__xnor2_1
XFILLER_87_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7016_ _7015_/A _7015_/C _7015_/B vssd1 vssd1 vccd1 vccd1 _7017_/C sky130_fd_sc_hd__a21o_1
XFILLER_28_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7918_ _8099_/B vssd1 vssd1 vccd1 vccd1 _7984_/C sky130_fd_sc_hd__clkbuf_2
X_7849_ _8317_/B _8147_/A vssd1 vssd1 vccd1 vccd1 _7855_/A sky130_fd_sc_hd__or2_1
XFILLER_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5200_ _8419_/A vssd1 vssd1 vccd1 vccd1 _5200_/X sky130_fd_sc_hd__clkbuf_2
X_6180_ _6163_/A _6178_/X _6179_/X vssd1 vssd1 vccd1 vccd1 _6182_/A sky130_fd_sc_hd__o21a_1
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5131_ _5131_/A _5131_/B _5131_/C vssd1 vssd1 vccd1 vccd1 _5131_/X sky130_fd_sc_hd__and3_1
XFILLER_69_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5062_ _5051_/A _5109_/C _5050_/X _5061_/X _5069_/A vssd1 vssd1 vccd1 vccd1 _5062_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_84_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8610__26 vssd1 vssd1 vccd1 vccd1 _8610__26/HI _8705_/A sky130_fd_sc_hd__conb_1
XFILLER_37_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8752_ _8752_/A _4353_/Y vssd1 vssd1 vccd1 vccd1 io_out[37] sky130_fd_sc_hd__ebufn_8
XFILLER_80_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5964_ _5961_/A _5961_/B _5963_/Y vssd1 vssd1 vccd1 vccd1 _5964_/Y sky130_fd_sc_hd__a21oi_1
X_7703_ _8370_/A _8370_/B vssd1 vssd1 vccd1 vccd1 _7707_/B sky130_fd_sc_hd__and2b_1
X_4915_ _4915_/A vssd1 vssd1 vccd1 vccd1 _5030_/B sky130_fd_sc_hd__buf_2
X_8683_ _8683_/A _4390_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[0] sky130_fd_sc_hd__ebufn_8
X_5895_ _5889_/A _5889_/B _5888_/A vssd1 vssd1 vccd1 vccd1 _5961_/A sky130_fd_sc_hd__o21ai_1
XFILLER_33_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4846_ _4873_/A vssd1 vssd1 vccd1 vccd1 _4848_/A sky130_fd_sc_hd__clkbuf_2
X_7634_ _7717_/B _7634_/B vssd1 vssd1 vccd1 vccd1 _7637_/A sky130_fd_sc_hd__xor2_1
X_7565_ _7733_/A vssd1 vssd1 vccd1 vccd1 _7620_/A sky130_fd_sc_hd__clkbuf_2
X_4777_ _4897_/A _4966_/A _4991_/A vssd1 vssd1 vccd1 vccd1 _4960_/A sky130_fd_sc_hd__or3_4
X_6516_ _8565_/Q vssd1 vssd1 vccd1 vccd1 _6521_/A sky130_fd_sc_hd__inv_2
XFILLER_20_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7496_ _7770_/A vssd1 vssd1 vccd1 vccd1 _7824_/A sky130_fd_sc_hd__clkbuf_2
X_6447_ _6442_/A _6442_/B _6440_/B vssd1 vssd1 vccd1 vccd1 _6448_/B sky130_fd_sc_hd__a21oi_1
X_6378_ _6380_/B _6380_/C _6326_/B vssd1 vssd1 vccd1 vccd1 _6378_/Y sky130_fd_sc_hd__o21ai_1
X_8117_ _8078_/A _8078_/B _8116_/X vssd1 vssd1 vccd1 vccd1 _8168_/A sky130_fd_sc_hd__a21oi_1
X_5329_ _8509_/Q vssd1 vssd1 vccd1 vccd1 _5374_/A sky130_fd_sc_hd__inv_2
X_8048_ _8048_/A _8048_/B vssd1 vssd1 vccd1 vccd1 _8048_/X sky130_fd_sc_hd__and2_1
XFILLER_87_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8676__92 vssd1 vssd1 vccd1 vccd1 _8676__92/HI _8785_/A sky130_fd_sc_hd__conb_1
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4700_ _4700_/A vssd1 vssd1 vccd1 vccd1 _8471_/D sky130_fd_sc_hd__clkbuf_1
X_5680_ _6082_/A _6248_/A _5591_/B _6090_/D vssd1 vssd1 vccd1 vccd1 _5681_/B sky130_fd_sc_hd__a31o_1
XFILLER_42_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4631_ _5441_/B _6482_/B _5121_/A vssd1 vssd1 vccd1 vccd1 _4950_/A sky130_fd_sc_hd__and3_1
XFILLER_8_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7350_ _7372_/A vssd1 vssd1 vccd1 vccd1 _7350_/Y sky130_fd_sc_hd__inv_2
X_4562_ _8448_/Q _4561_/B _4536_/X vssd1 vssd1 vccd1 vccd1 _4563_/B sky130_fd_sc_hd__o21ai_1
X_4493_ _8480_/Q _4495_/B vssd1 vssd1 vccd1 vccd1 _4494_/A sky130_fd_sc_hd__and2_1
X_7281_ _6912_/A _6912_/B _7280_/X vssd1 vssd1 vccd1 vccd1 _7334_/A sky130_fd_sc_hd__a21oi_1
X_6301_ _6301_/A _6301_/B vssd1 vssd1 vccd1 vccd1 _8526_/D sky130_fd_sc_hd__nor2_1
X_6232_ _6232_/A _6232_/B vssd1 vssd1 vccd1 vccd1 _6232_/Y sky130_fd_sc_hd__xnor2_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6163_ _6163_/A _6163_/B vssd1 vssd1 vccd1 vccd1 _6164_/B sky130_fd_sc_hd__xnor2_1
X_5114_ _5092_/C _5091_/X _5110_/X _4596_/A _5113_/X vssd1 vssd1 vccd1 vccd1 _5114_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_84_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6094_ _6069_/X _6232_/A _6232_/B _6093_/X vssd1 vssd1 vccd1 vccd1 _6241_/B sky130_fd_sc_hd__a31o_1
X_5045_ _5176_/S _5109_/B _5045_/C vssd1 vssd1 vccd1 vccd1 _5045_/X sky130_fd_sc_hd__or3_1
XFILLER_84_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6996_ _6996_/A _6996_/B _6996_/C vssd1 vssd1 vccd1 vccd1 _6996_/X sky130_fd_sc_hd__and3_1
XFILLER_53_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8735_ _8735_/A _4322_/Y vssd1 vssd1 vccd1 vccd1 io_out[20] sky130_fd_sc_hd__ebufn_8
XFILLER_53_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5947_ _5938_/A _5774_/A _5838_/A vssd1 vssd1 vccd1 vccd1 _6150_/A sky130_fd_sc_hd__a21o_1
X_5878_ _5984_/A vssd1 vssd1 vccd1 vccd1 _6184_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_21_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7617_ _7562_/A _7576_/A _7562_/C _7616_/Y vssd1 vssd1 vccd1 vccd1 _7618_/C sky130_fd_sc_hd__a31o_2
X_4829_ _4969_/B vssd1 vssd1 vccd1 vccd1 _5147_/B sky130_fd_sc_hd__clkbuf_2
X_7548_ _7549_/A _7549_/B _7547_/Y _7654_/B vssd1 vssd1 vccd1 vccd1 _7674_/A sky130_fd_sc_hd__a22oi_2
X_7479_ _8574_/Q _6348_/X _7478_/X vssd1 vssd1 vccd1 vccd1 _8574_/D sky130_fd_sc_hd__a21bo_1
XFILLER_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6850_ _6850_/A vssd1 vssd1 vccd1 vccd1 _7297_/A sky130_fd_sc_hd__clkbuf_4
X_6781_ _6781_/A _6781_/B vssd1 vssd1 vccd1 vccd1 _7279_/A sky130_fd_sc_hd__nand2_1
X_5801_ _5918_/C _5902_/A vssd1 vssd1 vccd1 vccd1 _5801_/Y sky130_fd_sc_hd__nand2_1
XFILLER_22_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5732_ _5825_/A _5824_/A vssd1 vssd1 vccd1 vccd1 _5733_/B sky130_fd_sc_hd__and2_1
X_8520_ input3/X _8520_/D vssd1 vssd1 vccd1 vccd1 _8520_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_50_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5663_ _5664_/A _5664_/B vssd1 vssd1 vccd1 vccd1 _5663_/Y sky130_fd_sc_hd__nor2_1
X_8451_ input3/X _8451_/D vssd1 vssd1 vccd1 vccd1 _8451_/Q sky130_fd_sc_hd__dfxtp_1
X_4614_ _4614_/A vssd1 vssd1 vccd1 vccd1 _5174_/S sky130_fd_sc_hd__clkbuf_2
X_8382_ _8384_/S _8381_/Y _8385_/A _8385_/B _8385_/C vssd1 vssd1 vccd1 vccd1 _8382_/X
+ sky130_fd_sc_hd__a2111o_1
X_5594_ _5664_/A vssd1 vssd1 vccd1 vccd1 _5594_/Y sky130_fd_sc_hd__inv_2
X_7402_ _7403_/A _7403_/B vssd1 vssd1 vccd1 vccd1 _7404_/A sky130_fd_sc_hd__nand2_1
X_7333_ _7333_/A _7333_/B vssd1 vssd1 vccd1 vccd1 _7334_/B sky130_fd_sc_hd__xnor2_1
X_4545_ _4548_/C _4545_/B vssd1 vssd1 vccd1 vccd1 _8442_/D sky130_fd_sc_hd__nor2_1
X_4476_ _8476_/Q _4480_/B vssd1 vssd1 vccd1 vccd1 _4477_/A sky130_fd_sc_hd__and2_1
X_7264_ _7264_/A _7264_/B _7264_/C vssd1 vssd1 vccd1 vccd1 _7265_/B sky130_fd_sc_hd__or3_1
X_7195_ _7196_/A _7196_/B _7196_/C vssd1 vssd1 vccd1 vccd1 _7200_/B sky130_fd_sc_hd__o21ai_2
X_6215_ _6215_/A _6215_/B vssd1 vssd1 vccd1 vccd1 _6222_/A sky130_fd_sc_hd__xnor2_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6146_ _6146_/A _6146_/B vssd1 vssd1 vccd1 vccd1 _6158_/A sky130_fd_sc_hd__xnor2_1
XINSDIODE2_25 _8708_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_14 _4445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_47 _8743_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6077_ _6088_/A _6088_/B vssd1 vssd1 vccd1 vccd1 _6079_/B sky130_fd_sc_hd__or2b_1
XINSDIODE2_58 _8775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_36 _8714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5028_ _8455_/Q _5030_/C _5041_/C _5028_/D vssd1 vssd1 vccd1 vccd1 _5028_/X sky130_fd_sc_hd__or4_1
XINSDIODE2_69 _8780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6979_ _6989_/A _6989_/B vssd1 vssd1 vccd1 vccd1 _7050_/A sky130_fd_sc_hd__xor2_2
XFILLER_13_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8718_ _8718_/A _4300_/Y vssd1 vssd1 vccd1 vccd1 io_out[3] sky130_fd_sc_hd__ebufn_8
XFILLER_70_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8646__62 vssd1 vssd1 vccd1 vccd1 _8646__62/HI _8755_/A sky130_fd_sc_hd__conb_1
XFILLER_88_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4330_ _4332_/A vssd1 vssd1 vccd1 vccd1 _4330_/Y sky130_fd_sc_hd__inv_2
X_4261_ _4264_/A vssd1 vssd1 vccd1 vccd1 _4261_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6000_ _6110_/B _6000_/B vssd1 vssd1 vccd1 vccd1 _6004_/A sky130_fd_sc_hd__nor2_1
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7951_ _7951_/A _8260_/A vssd1 vssd1 vccd1 vccd1 _7952_/C sky130_fd_sc_hd__nand2_1
X_6902_ _6930_/A _6902_/B vssd1 vssd1 vccd1 vccd1 _6904_/B sky130_fd_sc_hd__xnor2_2
X_7882_ _7880_/X _7856_/B _7881_/Y vssd1 vssd1 vccd1 vccd1 _7942_/A sky130_fd_sc_hd__a21bo_2
X_6833_ _6858_/A _6832_/C _6914_/B vssd1 vssd1 vccd1 vccd1 _6834_/C sky130_fd_sc_hd__a21o_1
XFILLER_23_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6764_ _6764_/A _6764_/B vssd1 vssd1 vccd1 vccd1 _6771_/A sky130_fd_sc_hd__xnor2_2
X_6695_ _6761_/A _6721_/B _6679_/B vssd1 vssd1 vccd1 vccd1 _6698_/B sky130_fd_sc_hd__o21ai_1
X_8503_ input3/X _8503_/D vssd1 vssd1 vccd1 vccd1 _8503_/Q sky130_fd_sc_hd__dfxtp_1
X_5715_ _5715_/A _5715_/B vssd1 vssd1 vccd1 vccd1 _5716_/B sky130_fd_sc_hd__or2_1
XFILLER_31_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5646_ _8515_/Q _7766_/B vssd1 vssd1 vccd1 vccd1 _5646_/Y sky130_fd_sc_hd__nor2_1
X_8434_ input3/X _8434_/D vssd1 vssd1 vccd1 vccd1 _8434_/Q sky130_fd_sc_hd__dfxtp_1
X_8365_ _8192_/X _8354_/Y _8363_/Y _8364_/X vssd1 vssd1 vccd1 vccd1 _8385_/C sky130_fd_sc_hd__a211o_2
X_5577_ _5577_/A _5679_/B vssd1 vssd1 vccd1 vccd1 _6082_/A sky130_fd_sc_hd__xnor2_2
X_7316_ _6795_/A _6794_/A _6794_/B _7315_/X vssd1 vssd1 vccd1 vccd1 _7318_/A sky130_fd_sc_hd__o31ai_1
X_8296_ _8286_/A _8296_/B vssd1 vssd1 vccd1 vccd1 _8298_/A sky130_fd_sc_hd__and2b_1
XFILLER_2_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4528_ _8437_/Q _4526_/A _4524_/X vssd1 vssd1 vccd1 vccd1 _4529_/B sky130_fd_sc_hd__o21ai_1
X_7247_ _7247_/A _7247_/B vssd1 vssd1 vccd1 vccd1 _7250_/B sky130_fd_sc_hd__and2_1
X_4459_ _5180_/B _4593_/A _4459_/C _4657_/A vssd1 vssd1 vccd1 vccd1 _4470_/B sky130_fd_sc_hd__or4_1
X_7178_ _7177_/A _7177_/B _7177_/C vssd1 vssd1 vccd1 vccd1 _7187_/B sky130_fd_sc_hd__a21o_1
X_6129_ _6129_/A _6129_/B vssd1 vssd1 vccd1 vccd1 _6130_/B sky130_fd_sc_hd__or2_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5500_ _5499_/A _5499_/C _5499_/B vssd1 vssd1 vccd1 vccd1 _5764_/C sky130_fd_sc_hd__a21oi_1
X_6480_ _6999_/A _6999_/B vssd1 vssd1 vccd1 vccd1 _6481_/A sky130_fd_sc_hd__xnor2_1
X_5431_ _8461_/Q _8524_/Q vssd1 vssd1 vccd1 vccd1 _5432_/B sky130_fd_sc_hd__or2b_1
X_8150_ _8258_/A _8258_/B vssd1 vssd1 vccd1 vccd1 _8152_/A sky130_fd_sc_hd__xnor2_1
X_5362_ _5362_/A _5367_/S _5362_/C _5366_/B vssd1 vssd1 vccd1 vccd1 _5363_/B sky130_fd_sc_hd__nand4_1
X_4313_ _4314_/A vssd1 vssd1 vccd1 vccd1 _4313_/Y sky130_fd_sc_hd__inv_2
X_7101_ _7101_/A _7040_/Y vssd1 vssd1 vccd1 vccd1 _7102_/B sky130_fd_sc_hd__or2b_1
X_8081_ _8084_/A _8084_/B vssd1 vssd1 vccd1 vccd1 _8082_/B sky130_fd_sc_hd__xor2_1
X_7032_ _7032_/A _7032_/B _7032_/C vssd1 vssd1 vccd1 vccd1 _7033_/B sky130_fd_sc_hd__nor3_1
X_5293_ _8505_/Q vssd1 vssd1 vccd1 vccd1 _5293_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7934_ _7934_/A _7934_/B vssd1 vssd1 vccd1 vccd1 _7935_/B sky130_fd_sc_hd__xor2_1
XFILLER_70_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7865_ _7865_/A _7865_/B vssd1 vssd1 vccd1 vccd1 _7866_/B sky130_fd_sc_hd__nand2_1
X_6816_ _6816_/A _6816_/B vssd1 vssd1 vccd1 vccd1 _6817_/C sky130_fd_sc_hd__nand2_1
XFILLER_23_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7796_ _7796_/A _7796_/B _7795_/Y vssd1 vssd1 vccd1 vccd1 _8213_/B sky130_fd_sc_hd__or3b_1
X_6747_ _6806_/A _7037_/A _6747_/C vssd1 vssd1 vccd1 vccd1 _6748_/B sky130_fd_sc_hd__and3b_1
XFILLER_50_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6678_ _6658_/A _6678_/B vssd1 vssd1 vccd1 vccd1 _6690_/A sky130_fd_sc_hd__and2b_1
X_5629_ _5754_/A _5629_/B vssd1 vssd1 vccd1 vccd1 _5631_/C sky130_fd_sc_hd__nand2_1
X_8417_ _8429_/S _8417_/B vssd1 vssd1 vccd1 vccd1 _8417_/X sky130_fd_sc_hd__and2_1
X_8348_ _8348_/A _8348_/B vssd1 vssd1 vccd1 vccd1 _8348_/X sky130_fd_sc_hd__xor2_2
X_8279_ _8279_/A _8279_/B vssd1 vssd1 vccd1 vccd1 _8334_/B sky130_fd_sc_hd__xnor2_1
X_8616__32 vssd1 vssd1 vccd1 vccd1 _8616__32/HI _8711_/A sky130_fd_sc_hd__conb_1
XFILLER_76_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5980_ _5918_/A _6106_/A _5980_/C vssd1 vssd1 vccd1 vccd1 _6106_/B sky130_fd_sc_hd__nand3b_1
XFILLER_37_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4931_ _5151_/A _4909_/B _4924_/X _4930_/X _4614_/A vssd1 vssd1 vccd1 vccd1 _4932_/C
+ sky130_fd_sc_hd__o311a_1
XFILLER_17_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4862_ _4862_/A _4862_/B vssd1 vssd1 vccd1 vccd1 _4863_/A sky130_fd_sc_hd__nor2_1
X_7650_ _7768_/A _8105_/A vssd1 vssd1 vccd1 vccd1 _7660_/A sky130_fd_sc_hd__nor2_1
XFILLER_60_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6601_ _7039_/B _6977_/B vssd1 vssd1 vccd1 vccd1 _6804_/B sky130_fd_sc_hd__nor2_1
XFILLER_20_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4793_ _4866_/A _5055_/B vssd1 vssd1 vccd1 vccd1 _5018_/A sky130_fd_sc_hd__or2_1
X_7581_ _7756_/A _7635_/C vssd1 vssd1 vccd1 vccd1 _7581_/Y sky130_fd_sc_hd__nor2_1
X_6532_ _7202_/A _6647_/A vssd1 vssd1 vccd1 vccd1 _6679_/B sky130_fd_sc_hd__or2_2
X_6463_ _6541_/A _7406_/A _6459_/Y _6461_/Y _6462_/X vssd1 vssd1 vccd1 vccd1 _8555_/D
+ sky130_fd_sc_hd__a221o_1
X_5414_ _5562_/A _5412_/B _5413_/X vssd1 vssd1 vccd1 vccd1 _5429_/A sky130_fd_sc_hd__a21bo_1
X_8202_ _8202_/A _8202_/B _8202_/C vssd1 vssd1 vccd1 vccd1 _8204_/A sky130_fd_sc_hd__nor3_1
X_6394_ _8503_/Q _8502_/Q _6393_/X vssd1 vssd1 vccd1 vccd1 _6399_/C sky130_fd_sc_hd__or3b_1
X_8133_ _8075_/A _8133_/B vssd1 vssd1 vccd1 vccd1 _8165_/A sky130_fd_sc_hd__and2b_1
X_5345_ _5359_/B _5345_/B vssd1 vssd1 vccd1 vccd1 _5347_/A sky130_fd_sc_hd__and2b_1
X_5276_ _5276_/A _5276_/B vssd1 vssd1 vccd1 vccd1 _8499_/D sky130_fd_sc_hd__nor2_1
X_8064_ _8064_/A _8064_/B vssd1 vssd1 vccd1 vccd1 _8136_/B sky130_fd_sc_hd__xor2_1
X_7015_ _7015_/A _7015_/B _7015_/C vssd1 vssd1 vccd1 vccd1 _7017_/B sky130_fd_sc_hd__nand3_4
XFILLER_68_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7917_ _7645_/B _7647_/B _7681_/B _7766_/Y vssd1 vssd1 vccd1 vccd1 _8099_/B sky130_fd_sc_hd__a211o_1
XFILLER_70_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7848_ _7881_/A _7881_/B vssd1 vssd1 vccd1 vccd1 _7856_/A sky130_fd_sc_hd__xnor2_1
X_7779_ _8176_/B _7779_/B vssd1 vssd1 vccd1 vccd1 _7780_/B sky130_fd_sc_hd__nor2_1
XFILLER_7_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5130_ _5048_/X _5128_/X _5130_/S vssd1 vssd1 vccd1 vccd1 _5131_/C sky130_fd_sc_hd__mux2_1
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5061_ _5135_/A _5054_/X _5057_/X _5132_/A _5060_/X vssd1 vssd1 vccd1 vccd1 _5061_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_57_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8751_ _8751_/A _4355_/Y vssd1 vssd1 vccd1 vccd1 io_out[36] sky130_fd_sc_hd__ebufn_8
XFILLER_52_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5963_ _5963_/A _5963_/B vssd1 vssd1 vccd1 vccd1 _5963_/Y sky130_fd_sc_hd__nor2_1
X_4914_ _4914_/A vssd1 vssd1 vccd1 vccd1 _4989_/A sky130_fd_sc_hd__clkbuf_2
X_7702_ _7702_/A _7702_/B vssd1 vssd1 vccd1 vccd1 _8370_/B sky130_fd_sc_hd__xor2_2
XFILLER_40_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5894_ _6065_/A _6065_/B vssd1 vssd1 vccd1 vccd1 _6067_/B sky130_fd_sc_hd__nor2_1
X_4845_ _5101_/S vssd1 vssd1 vccd1 vccd1 _4873_/A sky130_fd_sc_hd__buf_2
XFILLER_20_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7633_ _7633_/A _7633_/B vssd1 vssd1 vccd1 vccd1 _7634_/B sky130_fd_sc_hd__xnor2_1
X_4776_ _4805_/A _4908_/B vssd1 vssd1 vccd1 vccd1 _4991_/A sky130_fd_sc_hd__and2b_2
X_7564_ _8581_/Q _8457_/Q vssd1 vssd1 vccd1 vccd1 _7733_/A sky130_fd_sc_hd__xnor2_1
X_6515_ _6649_/B vssd1 vssd1 vccd1 vccd1 _6570_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_7495_ _7537_/A _7537_/B vssd1 vssd1 vccd1 vccd1 _7770_/A sky130_fd_sc_hd__and2_1
X_6446_ _6444_/Y _6446_/B vssd1 vssd1 vccd1 vccd1 _6448_/A sky130_fd_sc_hd__and2b_1
X_6377_ _6380_/C _6377_/B vssd1 vssd1 vccd1 vccd1 _8542_/D sky130_fd_sc_hd__nor2_1
X_5328_ _5328_/A vssd1 vssd1 vccd1 vccd1 _5333_/A sky130_fd_sc_hd__clkbuf_2
X_8116_ _8077_/A _8116_/B vssd1 vssd1 vccd1 vccd1 _8116_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8047_ _8047_/A _8047_/B vssd1 vssd1 vccd1 vccd1 _8078_/A sky130_fd_sc_hd__xor2_2
X_5259_ _6396_/D _5258_/C _8495_/Q vssd1 vssd1 vccd1 vccd1 _5261_/B sky130_fd_sc_hd__a21o_1
XFILLER_87_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4630_ _4623_/X _4629_/A _4629_/Y _4602_/X vssd1 vssd1 vccd1 vccd1 _8457_/D sky130_fd_sc_hd__o211a_1
XFILLER_30_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4561_ _8448_/Q _4561_/B vssd1 vssd1 vccd1 vccd1 _4566_/C sky130_fd_sc_hd__and2_1
X_6300_ _8526_/Q _5326_/B _6298_/X _6462_/A vssd1 vssd1 vccd1 vccd1 _6301_/B sky130_fd_sc_hd__a31o_1
X_7280_ _6911_/B _7280_/B vssd1 vssd1 vccd1 vccd1 _7280_/X sky130_fd_sc_hd__and2b_1
X_4492_ _4492_/A vssd1 vssd1 vccd1 vccd1 _8733_/A sky130_fd_sc_hd__clkbuf_1
X_6231_ _6232_/A _6232_/B _6081_/A vssd1 vssd1 vccd1 vccd1 _6231_/Y sky130_fd_sc_hd__a21oi_1
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6162_ _6162_/A _6179_/A vssd1 vssd1 vccd1 vccd1 _6163_/B sky130_fd_sc_hd__xnor2_1
X_5113_ _5113_/A _5113_/B vssd1 vssd1 vccd1 vccd1 _5113_/X sky130_fd_sc_hd__or2_1
XFILLER_69_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6093_ _6079_/A _6081_/A _6069_/B vssd1 vssd1 vccd1 vccd1 _6093_/X sky130_fd_sc_hd__o21a_1
X_5044_ _5080_/A _5034_/X _5043_/X _4863_/A vssd1 vssd1 vccd1 vccd1 _5045_/C sky130_fd_sc_hd__o211a_1
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6995_ _6996_/A _6996_/B _6996_/C vssd1 vssd1 vccd1 vccd1 _6995_/Y sky130_fd_sc_hd__a21oi_2
X_8734_ _8734_/A _4320_/Y vssd1 vssd1 vccd1 vccd1 io_out[19] sky130_fd_sc_hd__ebufn_8
X_5946_ _5833_/A _5833_/B _6154_/A vssd1 vssd1 vccd1 vccd1 _5952_/A sky130_fd_sc_hd__a21oi_1
X_5877_ _6118_/A _5899_/B vssd1 vssd1 vccd1 vccd1 _5880_/B sky130_fd_sc_hd__xor2_1
X_4828_ _5090_/A vssd1 vssd1 vccd1 vccd1 _5151_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_7616_ _7616_/A _7616_/B vssd1 vssd1 vccd1 vccd1 _7616_/Y sky130_fd_sc_hd__nand2_1
X_4759_ _4759_/A _4759_/B _4790_/B vssd1 vssd1 vccd1 vccd1 _4792_/A sky130_fd_sc_hd__or3_2
X_7547_ _7639_/A _7547_/B vssd1 vssd1 vccd1 vccd1 _7547_/Y sky130_fd_sc_hd__xnor2_1
X_7478_ _7478_/A _8430_/A _7478_/C _7488_/S vssd1 vssd1 vccd1 vccd1 _7478_/X sky130_fd_sc_hd__or4_1
X_6429_ _8550_/Q vssd1 vssd1 vccd1 vccd1 _6435_/A sky130_fd_sc_hd__inv_2
XFILLER_0_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6780_ _6780_/A _6781_/B vssd1 vssd1 vccd1 vccd1 _7328_/A sky130_fd_sc_hd__or2_1
X_5800_ _5800_/A _5800_/B vssd1 vssd1 vccd1 vccd1 _5902_/A sky130_fd_sc_hd__nand2_1
X_5731_ _5938_/A _5778_/A _6025_/B vssd1 vssd1 vccd1 vccd1 _5948_/A sky130_fd_sc_hd__nor3_2
X_8450_ input3/X _8450_/D vssd1 vssd1 vccd1 vccd1 _8450_/Q sky130_fd_sc_hd__dfxtp_1
X_5662_ _5662_/A _5662_/B vssd1 vssd1 vccd1 vccd1 _5667_/A sky130_fd_sc_hd__xnor2_1
XFILLER_30_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4613_ _4613_/A vssd1 vssd1 vccd1 vccd1 _8455_/D sky130_fd_sc_hd__clkbuf_1
X_7401_ _6521_/A _7403_/B _7409_/S vssd1 vssd1 vccd1 vccd1 _7405_/A sky130_fd_sc_hd__o21ai_1
X_8381_ _8381_/A _8381_/B vssd1 vssd1 vccd1 vccd1 _8381_/Y sky130_fd_sc_hd__nand2_1
X_5593_ _5593_/A vssd1 vssd1 vccd1 vccd1 _6259_/A sky130_fd_sc_hd__inv_2
X_7332_ _7332_/A _7332_/B vssd1 vssd1 vccd1 vccd1 _7333_/B sky130_fd_sc_hd__xnor2_1
X_4544_ _8442_/Q _4543_/B _4524_/X vssd1 vssd1 vccd1 vccd1 _4545_/B sky130_fd_sc_hd__o21ai_1
X_7263_ _7264_/A _7264_/B _7264_/C vssd1 vssd1 vccd1 vccd1 _7263_/X sky130_fd_sc_hd__o21a_1
X_4475_ _4475_/A vssd1 vssd1 vccd1 vccd1 _8729_/A sky130_fd_sc_hd__clkbuf_1
X_6214_ _6214_/A _6214_/B vssd1 vssd1 vccd1 vccd1 _6215_/B sky130_fd_sc_hd__xnor2_1
X_7194_ _7194_/A _7194_/B vssd1 vssd1 vccd1 vccd1 _7196_/C sky130_fd_sc_hd__xnor2_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6145_ _5932_/B _6021_/B _6020_/A vssd1 vssd1 vccd1 vccd1 _6146_/B sky130_fd_sc_hd__o21a_1
XINSDIODE2_15 _5055_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6076_ _6076_/A _6076_/B vssd1 vssd1 vccd1 vccd1 _6088_/B sky130_fd_sc_hd__xnor2_1
XINSDIODE2_37 _8714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5027_ _5148_/A _5104_/B _4906_/B _4848_/A vssd1 vssd1 vccd1 vccd1 _5027_/X sky130_fd_sc_hd__o31a_1
XINSDIODE2_59 _8775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_26 _8709_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_48 _8744_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8717_ _8717_/A _4299_/Y vssd1 vssd1 vccd1 vccd1 io_out[2] sky130_fd_sc_hd__ebufn_8
XFILLER_80_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6978_ _6978_/A _6978_/B vssd1 vssd1 vccd1 vccd1 _6989_/B sky130_fd_sc_hd__xnor2_2
XFILLER_13_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5929_ _6137_/B vssd1 vssd1 vccd1 vccd1 _5930_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_41_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8579_ input3/X _8579_/D vssd1 vssd1 vccd1 vccd1 _8579_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8661__77 vssd1 vssd1 vccd1 vccd1 _8661__77/HI _8770_/A sky130_fd_sc_hd__conb_1
XFILLER_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4260_ _4264_/A vssd1 vssd1 vccd1 vccd1 _4260_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7950_ _7950_/A vssd1 vssd1 vccd1 vccd1 _8053_/B sky130_fd_sc_hd__inv_2
XFILLER_82_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6901_ _6895_/Y _6924_/A _6900_/Y _6883_/X vssd1 vssd1 vccd1 vccd1 _6904_/A sky130_fd_sc_hd__a211oi_4
X_7881_ _7881_/A _7881_/B vssd1 vssd1 vccd1 vccd1 _7881_/Y sky130_fd_sc_hd__nand2_1
X_6832_ _6980_/A _6858_/A _6832_/C vssd1 vssd1 vccd1 vccd1 _6858_/B sky130_fd_sc_hd__nand3_1
XFILLER_35_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6763_ _6781_/A _6781_/B vssd1 vssd1 vccd1 vccd1 _6764_/B sky130_fd_sc_hd__xnor2_2
XFILLER_23_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6694_ _6694_/A vssd1 vssd1 vccd1 vccd1 _6721_/B sky130_fd_sc_hd__clkbuf_2
X_8502_ input3/X _8502_/D vssd1 vssd1 vccd1 vccd1 _8502_/Q sky130_fd_sc_hd__dfxtp_1
X_5714_ _5715_/A _5715_/B vssd1 vssd1 vccd1 vccd1 _5889_/A sky130_fd_sc_hd__nand2_1
X_5645_ _5686_/A _5684_/A vssd1 vssd1 vccd1 vccd1 _5659_/A sky130_fd_sc_hd__nand2_1
XFILLER_31_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8433_ input3/X _8433_/D vssd1 vssd1 vccd1 vccd1 _8433_/Q sky130_fd_sc_hd__dfxtp_1
X_8364_ _8364_/A _8364_/B vssd1 vssd1 vccd1 vccd1 _8364_/X sky130_fd_sc_hd__xor2_1
X_5576_ _5562_/A _5900_/A _5578_/B _5575_/A vssd1 vssd1 vccd1 vccd1 _5679_/B sky130_fd_sc_hd__a31o_1
X_7315_ _7315_/A _6798_/B vssd1 vssd1 vccd1 vccd1 _7315_/X sky130_fd_sc_hd__or2b_1
XFILLER_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8295_ _8295_/A _8290_/B vssd1 vssd1 vccd1 vccd1 _8300_/A sky130_fd_sc_hd__or2b_1
X_4527_ _8436_/Q _8437_/Q _4527_/C vssd1 vssd1 vccd1 vccd1 _4533_/C sky130_fd_sc_hd__and3_1
X_7246_ _7233_/A _7233_/B _7233_/C vssd1 vssd1 vccd1 vccd1 _7247_/B sky130_fd_sc_hd__o21ai_1
X_4458_ _4655_/A _6514_/A vssd1 vssd1 vccd1 vccd1 _4657_/A sky130_fd_sc_hd__or2_1
X_7177_ _7177_/A _7177_/B _7177_/C vssd1 vssd1 vccd1 vccd1 _7187_/A sky130_fd_sc_hd__nand3_1
X_4389_ _4390_/A vssd1 vssd1 vccd1 vccd1 _4389_/Y sky130_fd_sc_hd__inv_2
X_6128_ _6129_/A _6129_/B vssd1 vssd1 vccd1 vccd1 _6193_/A sky130_fd_sc_hd__nand2_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6059_ _6058_/A _6059_/B vssd1 vssd1 vccd1 vccd1 _6059_/X sky130_fd_sc_hd__and2b_1
XFILLER_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5430_ _8524_/Q _8461_/Q vssd1 vssd1 vccd1 vccd1 _5497_/A sky130_fd_sc_hd__or2b_1
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5361_ _5362_/A _5367_/S _5362_/C _5366_/B vssd1 vssd1 vccd1 vccd1 _5363_/A sky130_fd_sc_hd__a22o_1
X_4312_ _4314_/A vssd1 vssd1 vccd1 vccd1 _4312_/Y sky130_fd_sc_hd__inv_2
X_7100_ _7099_/A _7099_/B _7099_/C vssd1 vssd1 vccd1 vccd1 _7103_/B sky130_fd_sc_hd__a21o_1
X_5292_ _5292_/A vssd1 vssd1 vccd1 vccd1 _8504_/D sky130_fd_sc_hd__clkbuf_1
X_8080_ _8080_/A _8080_/B vssd1 vssd1 vccd1 vccd1 _8084_/B sky130_fd_sc_hd__xnor2_1
X_7031_ _6893_/A _6970_/B _6981_/S vssd1 vssd1 vccd1 vccd1 _7106_/A sky130_fd_sc_hd__o21ai_2
XFILLER_95_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7933_ _7933_/A _7933_/B vssd1 vssd1 vccd1 vccd1 _7934_/B sky130_fd_sc_hd__nand2_1
XFILLER_70_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7864_ _7864_/A _7864_/B _7864_/C vssd1 vssd1 vccd1 vccd1 _7865_/B sky130_fd_sc_hd__or3_1
X_6815_ _6839_/B _6814_/C _6814_/A vssd1 vssd1 vccd1 vccd1 _6817_/B sky130_fd_sc_hd__a21o_1
XFILLER_23_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7795_ _8193_/B _7795_/B vssd1 vssd1 vccd1 vccd1 _7795_/Y sky130_fd_sc_hd__nand2_1
X_6746_ _6751_/A _7033_/A vssd1 vssd1 vccd1 vccd1 _6747_/C sky130_fd_sc_hd__nand2_1
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6677_ _6678_/B _6669_/B _6676_/X vssd1 vssd1 vccd1 vccd1 _6777_/A sky130_fd_sc_hd__a21o_1
X_5628_ _5628_/A _5824_/A vssd1 vssd1 vccd1 vccd1 _5629_/B sky130_fd_sc_hd__nand2_1
X_8416_ _8415_/A _8415_/C _8415_/B vssd1 vssd1 vccd1 vccd1 _8417_/B sky130_fd_sc_hd__o21ai_1
X_8347_ _7983_/A _8249_/A _8306_/B _8041_/C vssd1 vssd1 vccd1 vccd1 _8348_/B sky130_fd_sc_hd__o22a_1
X_5559_ _5677_/B _5559_/B vssd1 vssd1 vccd1 vccd1 _5577_/A sky130_fd_sc_hd__or2_1
X_8278_ _8278_/A _8278_/B vssd1 vssd1 vccd1 vccd1 _8279_/B sky130_fd_sc_hd__or2_1
X_7229_ _7228_/B _7241_/A vssd1 vssd1 vccd1 vccd1 _7256_/B sky130_fd_sc_hd__and2b_1
XFILLER_86_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8631__47 vssd1 vssd1 vccd1 vccd1 _8631__47/HI _8740_/A sky130_fd_sc_hd__conb_1
XFILLER_61_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4930_ _5171_/A _4930_/B _5159_/B vssd1 vssd1 vccd1 vccd1 _4930_/X sky130_fd_sc_hd__or3_1
X_4861_ _4935_/A _4849_/X _4860_/X _5174_/S vssd1 vssd1 vccd1 vccd1 _4861_/X sky130_fd_sc_hd__o211a_1
XFILLER_17_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6600_ _7038_/B vssd1 vssd1 vccd1 vccd1 _6977_/B sky130_fd_sc_hd__clkbuf_2
X_4792_ _4792_/A _4798_/B vssd1 vssd1 vccd1 vccd1 _5055_/B sky130_fd_sc_hd__nor2_2
XFILLER_60_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7580_ _7725_/B vssd1 vssd1 vccd1 vccd1 _7635_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6531_ _6531_/A vssd1 vssd1 vccd1 vccd1 _6647_/A sky130_fd_sc_hd__buf_2
X_6462_ _6462_/A vssd1 vssd1 vccd1 vccd1 _6462_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_9_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6393_ _8501_/Q _8500_/Q _8505_/Q _8504_/Q vssd1 vssd1 vccd1 vccd1 _6393_/X sky130_fd_sc_hd__and4_1
X_5413_ _5565_/A _5565_/B vssd1 vssd1 vccd1 vccd1 _5413_/X sky130_fd_sc_hd__or2_1
X_8201_ _8201_/A _8201_/B _8201_/C vssd1 vssd1 vccd1 vccd1 _8202_/C sky130_fd_sc_hd__nor3_1
X_5344_ _5339_/B _5332_/X _5333_/X _5343_/Y vssd1 vssd1 vccd1 vccd1 _8511_/D sky130_fd_sc_hd__a22o_1
X_8132_ _8132_/A _8132_/B vssd1 vssd1 vccd1 vccd1 _8167_/A sky130_fd_sc_hd__nand2_1
X_5275_ _8499_/Q _5277_/C _5264_/X vssd1 vssd1 vccd1 vccd1 _5276_/B sky130_fd_sc_hd__o21ai_1
X_8063_ _8070_/A _8063_/B vssd1 vssd1 vccd1 vccd1 _8064_/B sky130_fd_sc_hd__xnor2_1
XFILLER_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7014_ _6948_/A _6947_/C _6947_/A vssd1 vssd1 vccd1 vccd1 _7015_/C sky130_fd_sc_hd__o21ai_2
XFILLER_68_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7916_ _7916_/A vssd1 vssd1 vccd1 vccd1 _8041_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_36_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7847_ _7886_/A _7847_/B vssd1 vssd1 vccd1 vccd1 _7881_/B sky130_fd_sc_hd__xnor2_1
XFILLER_23_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7778_ _7778_/A _7778_/B vssd1 vssd1 vccd1 vccd1 _7779_/B sky130_fd_sc_hd__and2_1
X_6729_ _6729_/A _6729_/B vssd1 vssd1 vccd1 vccd1 _6729_/Y sky130_fd_sc_hd__nor2_1
XFILLER_11_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5060_ _4596_/A _5087_/B _5080_/C _5058_/X _5059_/X vssd1 vssd1 vccd1 vccd1 _5060_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_96_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8750_ _8750_/A _4357_/Y vssd1 vssd1 vccd1 vccd1 io_out[35] sky130_fd_sc_hd__ebufn_8
XFILLER_65_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5962_ _6067_/A _6067_/B _6067_/C vssd1 vssd1 vccd1 vccd1 _6170_/A sky130_fd_sc_hd__o21a_1
X_4913_ _4913_/A vssd1 vssd1 vccd1 vccd1 _5104_/B sky130_fd_sc_hd__buf_2
XFILLER_18_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7701_ _8366_/A _8366_/B vssd1 vssd1 vccd1 vccd1 _8370_/A sky130_fd_sc_hd__or2_1
X_5893_ _5893_/A _5893_/B vssd1 vssd1 vccd1 vccd1 _6065_/B sky130_fd_sc_hd__xnor2_1
X_4844_ _5093_/A vssd1 vssd1 vccd1 vccd1 _5101_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_20_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7632_ _8367_/C _7756_/B _7632_/C vssd1 vssd1 vccd1 vccd1 _7633_/B sky130_fd_sc_hd__and3_1
X_4775_ _4944_/B _4804_/A vssd1 vssd1 vccd1 vccd1 _4966_/A sky130_fd_sc_hd__nor2_1
X_7563_ _7576_/A _7562_/C _7562_/A vssd1 vssd1 vccd1 vccd1 _7594_/B sky130_fd_sc_hd__a21o_1
X_6514_ _6514_/A _7403_/A vssd1 vssd1 vccd1 vccd1 _6649_/B sky130_fd_sc_hd__or2b_1
XFILLER_9_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7494_ _7494_/A _7494_/B vssd1 vssd1 vccd1 vccd1 _7537_/B sky130_fd_sc_hd__nand2_1
X_6445_ _6445_/A _6445_/B vssd1 vssd1 vccd1 vccd1 _6446_/B sky130_fd_sc_hd__nand2_1
X_6376_ _8542_/Q _6375_/B _6331_/B vssd1 vssd1 vccd1 vccd1 _6377_/B sky130_fd_sc_hd__o21ai_1
X_5327_ _6427_/A _5327_/B vssd1 vssd1 vccd1 vccd1 _5328_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8115_ _8115_/A _8115_/B vssd1 vssd1 vccd1 vccd1 _8169_/A sky130_fd_sc_hd__xnor2_1
X_8046_ _8046_/A _8046_/B vssd1 vssd1 vccd1 vccd1 _8047_/B sky130_fd_sc_hd__xnor2_2
XFILLER_87_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5258_ _8495_/Q _8494_/Q _5258_/C vssd1 vssd1 vccd1 vccd1 _5263_/B sky130_fd_sc_hd__and3_1
X_5189_ _8474_/Q _5192_/B vssd1 vssd1 vccd1 vccd1 _5189_/X sky130_fd_sc_hd__or2_1
XFILLER_28_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8601__17 vssd1 vssd1 vccd1 vccd1 _8601__17/HI _8696_/A sky130_fd_sc_hd__conb_1
XFILLER_83_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4560_ _4560_/A vssd1 vssd1 vccd1 vccd1 _8447_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4491_ _8479_/Q _4491_/B vssd1 vssd1 vccd1 vccd1 _4492_/A sky130_fd_sc_hd__and2_1
XFILLER_6_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6230_ _6230_/A _6230_/B vssd1 vssd1 vccd1 vccd1 _6264_/B sky130_fd_sc_hd__xnor2_4
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6161_ _6040_/A _6159_/X _6160_/X vssd1 vssd1 vccd1 vccd1 _6179_/A sky130_fd_sc_hd__o21a_1
X_8667__83 vssd1 vssd1 vccd1 vccd1 _8667__83/HI _8776_/A sky130_fd_sc_hd__conb_1
X_5112_ _5112_/A _5112_/B _5156_/B _5112_/D vssd1 vssd1 vccd1 vccd1 _5113_/B sky130_fd_sc_hd__or4_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6092_ _6238_/A _6238_/B _6089_/X _6091_/X vssd1 vssd1 vccd1 vccd1 _6232_/B sky130_fd_sc_hd__a31o_1
X_5043_ _5038_/X _5042_/X _5050_/A _5117_/B vssd1 vssd1 vccd1 vccd1 _5043_/X sky130_fd_sc_hd__a211o_1
XFILLER_84_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6994_ _7062_/A _7062_/B vssd1 vssd1 vccd1 vccd1 _6994_/Y sky130_fd_sc_hd__nand2_2
XFILLER_80_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8733_ _8733_/A _4319_/Y vssd1 vssd1 vccd1 vccd1 io_out[18] sky130_fd_sc_hd__ebufn_8
X_5945_ _5945_/A _5945_/B vssd1 vssd1 vccd1 vccd1 _5953_/A sky130_fd_sc_hd__xnor2_2
X_5876_ _5689_/A _6126_/A _5875_/X vssd1 vssd1 vccd1 vccd1 _5899_/B sky130_fd_sc_hd__o21ai_1
XFILLER_21_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4827_ _5138_/A _5138_/B _5138_/C _4609_/A vssd1 vssd1 vccd1 vccd1 _4827_/X sky130_fd_sc_hd__o31a_1
X_7615_ _7613_/X _7615_/B vssd1 vssd1 vccd1 vccd1 _7618_/B sky130_fd_sc_hd__and2b_1
XFILLER_21_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4758_ _4675_/B _4762_/A _4759_/B vssd1 vssd1 vccd1 vccd1 _4812_/A sky130_fd_sc_hd__and3b_1
XFILLER_5_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7546_ _7546_/A _7546_/B vssd1 vssd1 vccd1 vccd1 _7547_/B sky130_fd_sc_hd__xnor2_1
X_4689_ _4689_/A vssd1 vssd1 vccd1 vccd1 _7412_/A sky130_fd_sc_hd__clkbuf_2
X_7477_ _7477_/A _7477_/B _7477_/C vssd1 vssd1 vccd1 vccd1 _7488_/S sky130_fd_sc_hd__and3_1
XFILLER_4_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6428_ _6428_/A vssd1 vssd1 vccd1 vccd1 _6432_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6359_ _6362_/C _6359_/B vssd1 vssd1 vccd1 vccd1 _8536_/D sky130_fd_sc_hd__nor2_1
XFILLER_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8029_ _7984_/A _7983_/B _7982_/B _7986_/A _7986_/B vssd1 vssd1 vccd1 vccd1 _8091_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_84_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5730_ _5767_/B vssd1 vssd1 vccd1 vccd1 _6025_/B sky130_fd_sc_hd__clkbuf_2
X_7400_ _6432_/A _7409_/S _7398_/Y _7399_/X vssd1 vssd1 vccd1 vccd1 _8565_/D sky130_fd_sc_hd__a31o_1
X_5661_ _5685_/C _5661_/B vssd1 vssd1 vccd1 vccd1 _5662_/B sky130_fd_sc_hd__xnor2_1
X_4612_ _4657_/B _4612_/B _4643_/A vssd1 vssd1 vccd1 vccd1 _4613_/A sky130_fd_sc_hd__and3_1
X_8380_ _8381_/A _8381_/B vssd1 vssd1 vccd1 vccd1 _8384_/S sky130_fd_sc_hd__or2_1
X_5592_ _6082_/B _5592_/B vssd1 vssd1 vccd1 vccd1 _5593_/A sky130_fd_sc_hd__nor2_1
X_7331_ _7331_/A _7331_/B vssd1 vssd1 vccd1 vccd1 _7332_/B sky130_fd_sc_hd__xnor2_1
X_4543_ _8442_/Q _4543_/B vssd1 vssd1 vccd1 vccd1 _4548_/C sky130_fd_sc_hd__and2_1
X_7262_ _7146_/A _7146_/C _7146_/B vssd1 vssd1 vccd1 vccd1 _7264_/C sky130_fd_sc_hd__a21boi_1
X_4474_ _8475_/Q _4480_/B vssd1 vssd1 vccd1 vccd1 _4475_/A sky130_fd_sc_hd__and2_1
X_6213_ _6213_/A _6213_/B vssd1 vssd1 vccd1 vccd1 _6214_/B sky130_fd_sc_hd__xnor2_1
X_7193_ _7193_/A _7193_/B vssd1 vssd1 vccd1 vccd1 _7194_/A sky130_fd_sc_hd__nand2_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6144_ _6144_/A _6144_/B vssd1 vssd1 vccd1 vccd1 _6146_/A sky130_fd_sc_hd__nand2_1
XFILLER_57_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6075_ _6075_/A _6075_/B vssd1 vssd1 vccd1 vccd1 _6076_/A sky130_fd_sc_hd__nand2_1
XINSDIODE2_16 _8704_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_49 _8744_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_27 _8709_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5026_ _5026_/A vssd1 vssd1 vccd1 vccd1 _5148_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_57_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_38 _8715_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6977_ _6977_/A _6977_/B vssd1 vssd1 vccd1 vccd1 _6978_/B sky130_fd_sc_hd__nor2_1
X_8716_ _8716_/A _4298_/Y vssd1 vssd1 vccd1 vccd1 io_out[1] sky130_fd_sc_hd__ebufn_8
X_5928_ _5843_/A _5843_/B _5927_/X vssd1 vssd1 vccd1 vccd1 _5935_/A sky130_fd_sc_hd__a21bo_1
XFILLER_80_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5859_ _5918_/C _5859_/B vssd1 vssd1 vccd1 vccd1 _5863_/A sky130_fd_sc_hd__xor2_1
X_8578_ input3/X _8578_/D vssd1 vssd1 vccd1 vccd1 _8578_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_5_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7529_ _7655_/A _7654_/B vssd1 vssd1 vccd1 vccd1 _7682_/A sky130_fd_sc_hd__or2_1
XFILLER_79_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8637__53 vssd1 vssd1 vccd1 vccd1 _8637__53/HI _8746_/A sky130_fd_sc_hd__conb_1
XFILLER_67_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6900_ _6883_/A _6883_/C _6883_/D _6883_/B vssd1 vssd1 vccd1 vccd1 _6900_/Y sky130_fd_sc_hd__a22oi_4
X_7880_ _7881_/A _7881_/B vssd1 vssd1 vccd1 vccd1 _7880_/X sky130_fd_sc_hd__or2_1
X_6831_ _6874_/A _6831_/B vssd1 vssd1 vccd1 vccd1 _6838_/A sky130_fd_sc_hd__xor2_2
XFILLER_35_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8501_ input3/X _8501_/D vssd1 vssd1 vccd1 vccd1 _8501_/Q sky130_fd_sc_hd__dfxtp_1
X_6762_ _7026_/A _6778_/B vssd1 vssd1 vccd1 vccd1 _6764_/A sky130_fd_sc_hd__xnor2_2
XFILLER_50_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6693_ _6714_/B _6714_/C _6693_/C vssd1 vssd1 vccd1 vccd1 _6694_/A sky130_fd_sc_hd__or3_1
XFILLER_50_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5713_ _5914_/A _5713_/B vssd1 vssd1 vccd1 vccd1 _5715_/B sky130_fd_sc_hd__nor2_1
X_5644_ _5579_/B _5643_/Y _5535_/B _5541_/B vssd1 vssd1 vccd1 vccd1 _5683_/A sky130_fd_sc_hd__a22o_1
X_8432_ _7416_/X _8430_/Y _8431_/Y vssd1 vssd1 vccd1 vccd1 _8587_/D sky130_fd_sc_hd__a21oi_1
X_8363_ _8192_/X _8354_/Y _8355_/Y _8358_/Y _8362_/X vssd1 vssd1 vccd1 vccd1 _8363_/Y
+ sky130_fd_sc_hd__o2111ai_1
X_7314_ _7314_/A _7314_/B vssd1 vssd1 vccd1 vccd1 _7333_/A sky130_fd_sc_hd__xnor2_1
X_5575_ _5575_/A _5575_/B vssd1 vssd1 vccd1 vccd1 _5578_/B sky130_fd_sc_hd__nor2_1
X_4526_ _4526_/A _4526_/B vssd1 vssd1 vccd1 vccd1 _8436_/D sky130_fd_sc_hd__nor2_1
X_8294_ _8364_/A _8364_/B _8359_/C _8293_/Y _8291_/B vssd1 vssd1 vccd1 vccd1 _8353_/A
+ sky130_fd_sc_hd__a32o_2
X_7245_ _7253_/A _7253_/B vssd1 vssd1 vccd1 vccd1 _7351_/A sky130_fd_sc_hd__nor2_1
X_4457_ _4624_/A _4614_/A _5132_/A _4949_/A vssd1 vssd1 vccd1 vccd1 _4459_/C sky130_fd_sc_hd__o31a_1
X_7176_ _7176_/A _7176_/B _7206_/B vssd1 vssd1 vccd1 vccd1 _7177_/C sky130_fd_sc_hd__and3_1
X_4388_ _4390_/A vssd1 vssd1 vccd1 vccd1 _4388_/Y sky130_fd_sc_hd__inv_2
X_6127_ _5860_/B _6184_/B _6104_/Y vssd1 vssd1 vccd1 vccd1 _6129_/B sky130_fd_sc_hd__o21a_1
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6058_ _6058_/A _6059_/B vssd1 vssd1 vccd1 vccd1 _6071_/B sky130_fd_sc_hd__xnor2_1
X_5009_ _5050_/A _5058_/B _5009_/C _5009_/D vssd1 vssd1 vccd1 vccd1 _5009_/X sky130_fd_sc_hd__or4_1
XFILLER_38_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5360_ _5360_/A _5360_/B vssd1 vssd1 vccd1 vccd1 _5366_/B sky130_fd_sc_hd__or2_1
X_4311_ _4314_/A vssd1 vssd1 vccd1 vccd1 _4311_/Y sky130_fd_sc_hd__inv_2
X_5291_ _5291_/A _5291_/B _5291_/C vssd1 vssd1 vccd1 vccd1 _5292_/A sky130_fd_sc_hd__and3_1
X_7030_ _7272_/A _7030_/B vssd1 vssd1 vccd1 vccd1 _7030_/X sky130_fd_sc_hd__xor2_1
XFILLER_4_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7932_ _7932_/A _7932_/B vssd1 vssd1 vccd1 vccd1 _7933_/A sky130_fd_sc_hd__nand2_1
XFILLER_70_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7863_ _7864_/A _7864_/B _7864_/C vssd1 vssd1 vccd1 vccd1 _7865_/A sky130_fd_sc_hd__o21ai_1
XFILLER_35_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6814_ _6814_/A _6839_/B _6814_/C vssd1 vssd1 vccd1 vccd1 _6826_/A sky130_fd_sc_hd__nand3_1
X_7794_ _7796_/A _7796_/B _8193_/B _7795_/B vssd1 vssd1 vccd1 vccd1 _8210_/A sky130_fd_sc_hd__o211a_1
X_6745_ _6914_/A _6745_/B vssd1 vssd1 vccd1 vccd1 _7037_/A sky130_fd_sc_hd__nand2_1
XFILLER_50_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6676_ _6703_/B _6703_/A vssd1 vssd1 vccd1 vccd1 _6676_/X sky130_fd_sc_hd__and2b_1
X_8415_ _8415_/A _8415_/B _8415_/C vssd1 vssd1 vccd1 vccd1 _8429_/S sky130_fd_sc_hd__or3_1
X_5627_ _5627_/A vssd1 vssd1 vccd1 vccd1 _5824_/A sky130_fd_sc_hd__clkbuf_2
X_8346_ _8346_/A _8289_/B vssd1 vssd1 vccd1 vccd1 _8346_/X sky130_fd_sc_hd__or2b_1
X_5558_ _5677_/A _5557_/C _5557_/A vssd1 vssd1 vccd1 vccd1 _5559_/B sky130_fd_sc_hd__o21a_1
X_4509_ _5327_/B vssd1 vssd1 vccd1 vccd1 _5368_/B sky130_fd_sc_hd__clkbuf_2
X_8277_ _8277_/A _8277_/B vssd1 vssd1 vccd1 vccd1 _8278_/B sky130_fd_sc_hd__and2_1
XFILLER_2_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7228_ _7228_/A _7228_/B _7228_/C vssd1 vssd1 vccd1 vccd1 _7241_/A sky130_fd_sc_hd__or3_1
XFILLER_78_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5489_ _5487_/X _5488_/Y _5615_/A vssd1 vssd1 vccd1 vccd1 _5490_/B sky130_fd_sc_hd__mux2_1
XFILLER_76_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7159_ _7177_/A _7159_/B vssd1 vssd1 vccd1 vccd1 _7159_/X sky130_fd_sc_hd__and2b_1
XFILLER_46_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8607__23 vssd1 vssd1 vccd1 vccd1 _8607__23/HI _8702_/A sky130_fd_sc_hd__conb_1
XFILLER_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4860_ _4592_/A _5135_/C _4859_/X _4609_/A vssd1 vssd1 vccd1 vccd1 _4860_/X sky130_fd_sc_hd__a211o_1
XFILLER_32_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4791_ _4791_/A _4818_/B vssd1 vssd1 vccd1 vccd1 _4866_/A sky130_fd_sc_hd__nor2_1
X_6530_ _6761_/A vssd1 vssd1 vccd1 vccd1 _6721_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_60_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6461_ _7406_/A _6461_/B vssd1 vssd1 vccd1 vccd1 _6461_/Y sky130_fd_sc_hd__nor2_1
X_6392_ _8493_/Q _8492_/Q _6392_/C _8496_/Q vssd1 vssd1 vccd1 vccd1 _6399_/B sky130_fd_sc_hd__nand4_1
X_5412_ _5562_/A _5412_/B vssd1 vssd1 vccd1 vccd1 _5565_/B sky130_fd_sc_hd__xnor2_1
X_8200_ _8211_/A _8211_/B vssd1 vssd1 vccd1 vccd1 _8202_/B sky130_fd_sc_hd__or2b_1
X_5343_ _5343_/A _5343_/B vssd1 vssd1 vccd1 vccd1 _5343_/Y sky130_fd_sc_hd__xnor2_1
X_8131_ _8131_/A _8131_/B vssd1 vssd1 vccd1 vccd1 _8132_/B sky130_fd_sc_hd__or2_1
XFILLER_87_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5274_ _8499_/Q _5277_/C vssd1 vssd1 vccd1 vccd1 _5276_/A sky130_fd_sc_hd__and2_1
X_8062_ _7621_/B _8063_/B _7947_/X _8326_/A vssd1 vssd1 vccd1 vccd1 _8136_/A sky130_fd_sc_hd__o22ai_2
X_7013_ _7058_/A _7131_/A _6993_/B _6992_/B _6992_/A vssd1 vssd1 vccd1 vccd1 _7015_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_83_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7915_ _7915_/A _8299_/A vssd1 vssd1 vccd1 vccd1 _7930_/C sky130_fd_sc_hd__xnor2_1
X_7846_ _7860_/A _7844_/Y _7845_/X vssd1 vssd1 vccd1 vccd1 _7847_/B sky130_fd_sc_hd__a21o_1
X_4989_ _4989_/A _5009_/C vssd1 vssd1 vccd1 vccd1 _5004_/C sky130_fd_sc_hd__or2_1
XFILLER_11_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7777_ _7778_/A _7778_/B vssd1 vssd1 vccd1 vccd1 _8176_/B sky130_fd_sc_hd__nor2_1
X_6728_ _6729_/A _6729_/B vssd1 vssd1 vccd1 vccd1 _6951_/B sky130_fd_sc_hd__xnor2_1
X_6659_ _6660_/A _6660_/B vssd1 vssd1 vccd1 vccd1 _6886_/A sky130_fd_sc_hd__nand2_1
X_8329_ _8329_/A _8329_/B vssd1 vssd1 vccd1 vccd1 _8329_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_3_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5961_ _5961_/A _5961_/B vssd1 vssd1 vccd1 vccd1 _6067_/C sky130_fd_sc_hd__xor2_1
XFILLER_18_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4912_ _5135_/B _4907_/X _4975_/C _4911_/X _5179_/A vssd1 vssd1 vccd1 vccd1 _4932_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_52_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7700_ _8052_/A _8052_/B vssd1 vssd1 vccd1 vccd1 _8366_/B sky130_fd_sc_hd__or2_1
X_7631_ _8146_/A _8146_/B _8326_/A vssd1 vssd1 vccd1 vccd1 _7632_/C sky130_fd_sc_hd__o21ai_2
X_5892_ _5892_/A _5892_/B _5748_/B vssd1 vssd1 vccd1 vccd1 _6065_/A sky130_fd_sc_hd__or3b_1
X_4843_ _8454_/Q vssd1 vssd1 vccd1 vccd1 _5093_/A sky130_fd_sc_hd__inv_2
XFILLER_21_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4774_ _4786_/B vssd1 vssd1 vccd1 vccd1 _4944_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_60_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7562_ _7562_/A _7576_/A _7562_/C vssd1 vssd1 vccd1 vccd1 _7594_/A sky130_fd_sc_hd__nand3_1
X_6513_ _6570_/A vssd1 vssd1 vccd1 vccd1 _6513_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7493_ _7493_/A vssd1 vssd1 vccd1 vccd1 _7537_/A sky130_fd_sc_hd__buf_2
X_6444_ _6445_/A _6450_/B vssd1 vssd1 vccd1 vccd1 _6444_/Y sky130_fd_sc_hd__nor2_1
XFILLER_9_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6375_ _8542_/Q _6375_/B vssd1 vssd1 vccd1 vccd1 _6380_/C sky130_fd_sc_hd__and2_1
X_5326_ _7478_/A _5326_/B vssd1 vssd1 vccd1 vccd1 _5332_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8114_ _8114_/A _8114_/B vssd1 vssd1 vccd1 vccd1 _8115_/B sky130_fd_sc_hd__xor2_2
X_5257_ _6396_/D _5258_/C _5256_/Y vssd1 vssd1 vccd1 vccd1 _8494_/D sky130_fd_sc_hd__a21oi_1
X_8045_ _8131_/A _8045_/B vssd1 vssd1 vccd1 vccd1 _8046_/B sky130_fd_sc_hd__nor2_2
X_5188_ _5202_/A vssd1 vssd1 vccd1 vccd1 _5188_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_68_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8598__14 vssd1 vssd1 vccd1 vccd1 _8598__14/HI _8693_/A sky130_fd_sc_hd__conb_1
XFILLER_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7829_ _7926_/A _7830_/B _7826_/Y _7827_/X _7984_/A vssd1 vssd1 vccd1 vccd1 _8037_/A
+ sky130_fd_sc_hd__o2111a_1
XFILLER_22_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4490_ _4490_/A vssd1 vssd1 vccd1 vccd1 _8732_/A sky130_fd_sc_hd__clkbuf_1
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6160_ _6160_/A _6160_/B vssd1 vssd1 vccd1 vccd1 _6160_/X sky130_fd_sc_hd__or2_1
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5111_ _5148_/C _5092_/D _5014_/D vssd1 vssd1 vccd1 vccd1 _5113_/A sky130_fd_sc_hd__o21a_1
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6091_ _6233_/A _6090_/X _6233_/B vssd1 vssd1 vccd1 vccd1 _6091_/X sky130_fd_sc_hd__o21ba_1
X_8682__98 vssd1 vssd1 vccd1 vccd1 _8682__98/HI _8506_/D sky130_fd_sc_hd__conb_1
X_5042_ _4973_/A _5117_/C _5118_/A _5041_/X _4939_/X vssd1 vssd1 vccd1 vccd1 _5042_/X
+ sky130_fd_sc_hd__a2111o_1
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6993_ _6993_/A _6993_/B vssd1 vssd1 vccd1 vccd1 _7062_/B sky130_fd_sc_hd__xnor2_1
X_8732_ _8732_/A _4318_/Y vssd1 vssd1 vccd1 vccd1 io_out[17] sky130_fd_sc_hd__ebufn_8
X_5944_ _6015_/A _6015_/B vssd1 vssd1 vccd1 vccd1 _5945_/B sky130_fd_sc_hd__xnor2_1
XFILLER_43_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5875_ _5918_/A _5803_/B vssd1 vssd1 vccd1 vccd1 _5875_/X sky130_fd_sc_hd__or2b_1
X_4826_ _5132_/B _5051_/A vssd1 vssd1 vccd1 vccd1 _5138_/C sky130_fd_sc_hd__or2_1
X_7614_ _8463_/Q _8587_/Q vssd1 vssd1 vccd1 vccd1 _7615_/B sky130_fd_sc_hd__or2b_2
X_7545_ _7768_/A _7978_/A vssd1 vssd1 vccd1 vccd1 _7546_/B sky130_fd_sc_hd__nor2_1
X_4757_ _4908_/A _4749_/A _4908_/B vssd1 vssd1 vccd1 vccd1 _4772_/A sky130_fd_sc_hd__o21a_1
X_4688_ _7501_/B _4690_/B vssd1 vssd1 vccd1 vccd1 _4698_/C sky130_fd_sc_hd__nor2_1
X_7476_ _7477_/A _7477_/B _7477_/C vssd1 vssd1 vccd1 vccd1 _7478_/C sky130_fd_sc_hd__a21oi_1
X_6427_ _6427_/A _6465_/A vssd1 vssd1 vccd1 vccd1 _6428_/A sky130_fd_sc_hd__nor2_1
X_6358_ _8536_/Q _6356_/A _6331_/B vssd1 vssd1 vccd1 vccd1 _6359_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5309_ _5495_/A _5322_/C _6293_/B vssd1 vssd1 vccd1 vccd1 _5309_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_88_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6289_ _6289_/A _6289_/B _6289_/C _6289_/D vssd1 vssd1 vccd1 vccd1 _6298_/S sky130_fd_sc_hd__or4_1
X_8028_ _8341_/A _8028_/B vssd1 vssd1 vccd1 vccd1 _8091_/A sky130_fd_sc_hd__xnor2_1
XFILLER_29_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5660_ _6053_/B _5660_/B vssd1 vssd1 vccd1 vccd1 _5661_/B sky130_fd_sc_hd__nor2_1
XFILLER_30_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4611_ _4619_/A _4619_/B vssd1 vssd1 vccd1 vccd1 _4643_/A sky130_fd_sc_hd__or2_1
X_5591_ _6248_/A _5591_/B vssd1 vssd1 vccd1 vccd1 _5592_/B sky130_fd_sc_hd__nor2_1
XFILLER_30_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7330_ _7330_/A _7330_/B vssd1 vssd1 vccd1 vccd1 _7331_/B sky130_fd_sc_hd__xnor2_1
X_4542_ _4542_/A vssd1 vssd1 vccd1 vccd1 _8441_/D sky130_fd_sc_hd__clkbuf_1
X_7261_ _7098_/B _7093_/C _7093_/A vssd1 vssd1 vccd1 vccd1 _7264_/B sky130_fd_sc_hd__o21a_1
X_4473_ _4473_/A vssd1 vssd1 vccd1 vccd1 _8728_/A sky130_fd_sc_hd__clkbuf_1
X_6212_ _6114_/A _6114_/B _6211_/Y vssd1 vssd1 vccd1 vccd1 _6213_/B sky130_fd_sc_hd__a21bo_1
X_7192_ _7212_/A _7212_/B vssd1 vssd1 vccd1 vccd1 _7196_/B sky130_fd_sc_hd__and2_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6143_ _6143_/A _6143_/B vssd1 vssd1 vccd1 vccd1 _6144_/B sky130_fd_sc_hd__or2_1
XFILLER_85_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6074_ _6084_/A _6084_/B _6073_/X vssd1 vssd1 vccd1 vccd1 _6088_/A sky130_fd_sc_hd__o21a_1
X_8593__9 vssd1 vssd1 vccd1 vccd1 _8593__9/HI _8688_/A sky130_fd_sc_hd__conb_1
XINSDIODE2_39 _8715_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5025_ _5025_/A vssd1 vssd1 vccd1 vccd1 _5109_/C sky130_fd_sc_hd__clkbuf_2
XINSDIODE2_17 _8704_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_28 _8710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6976_ _6967_/X _7035_/B _6975_/X vssd1 vssd1 vccd1 vccd1 _6989_/A sky130_fd_sc_hd__a21oi_2
XFILLER_26_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8715_ _8715_/A _4388_/Y vssd1 vssd1 vccd1 vccd1 io_out[0] sky130_fd_sc_hd__ebufn_8
XFILLER_53_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5927_ _5927_/A _5842_/B vssd1 vssd1 vccd1 vccd1 _5927_/X sky130_fd_sc_hd__or2b_1
XFILLER_41_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5858_ _5694_/A _5804_/B _5999_/A _5857_/Y vssd1 vssd1 vccd1 vccd1 _5859_/B sky130_fd_sc_hd__a31o_1
XFILLER_21_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4809_ _4817_/A _4809_/B vssd1 vssd1 vccd1 vccd1 _4969_/A sky130_fd_sc_hd__nor2_1
X_8577_ input3/X _8577_/D vssd1 vssd1 vccd1 vccd1 _8577_/Q sky130_fd_sc_hd__dfxtp_1
X_5789_ _5818_/A _5818_/B vssd1 vssd1 vccd1 vccd1 _5814_/A sky130_fd_sc_hd__xnor2_1
X_7528_ _7813_/A _7528_/B _7528_/C vssd1 vssd1 vccd1 vccd1 _7654_/B sky130_fd_sc_hd__and3_1
X_7459_ _7459_/A _7459_/B vssd1 vssd1 vccd1 vccd1 _7461_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8652__68 vssd1 vssd1 vccd1 vccd1 _8652__68/HI _8761_/A sky130_fd_sc_hd__conb_1
XFILLER_82_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6830_ _6735_/Y _6736_/X _6858_/A _6832_/C vssd1 vssd1 vccd1 vccd1 _6831_/B sky130_fd_sc_hd__a22o_1
XFILLER_90_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6761_ _6761_/A _6780_/A vssd1 vssd1 vccd1 vccd1 _6778_/B sky130_fd_sc_hd__xnor2_2
XFILLER_90_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8500_ input3/X _8500_/D vssd1 vssd1 vccd1 vccd1 _8500_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5712_ _5707_/Y _5708_/X _5711_/Y _5860_/A vssd1 vssd1 vccd1 vccd1 _5713_/B sky130_fd_sc_hd__o2bb2a_1
X_6692_ _6777_/A _6777_/B vssd1 vssd1 vccd1 vccd1 _6796_/A sky130_fd_sc_hd__xnor2_1
XFILLER_31_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5643_ _5705_/A _5976_/A vssd1 vssd1 vccd1 vccd1 _5643_/Y sky130_fd_sc_hd__nor2_1
X_8431_ _7416_/X _8430_/Y _4510_/A vssd1 vssd1 vccd1 vccd1 _8431_/Y sky130_fd_sc_hd__o21ai_1
X_8362_ _8362_/A _8362_/B _8362_/C vssd1 vssd1 vccd1 vccd1 _8362_/X sky130_fd_sc_hd__and3_1
X_5574_ _5574_/A _5574_/B vssd1 vssd1 vccd1 vccd1 _5575_/B sky130_fd_sc_hd__and2_1
X_7313_ _7313_/A _7313_/B vssd1 vssd1 vccd1 vccd1 _7314_/B sky130_fd_sc_hd__xnor2_1
X_4525_ _8436_/Q _4527_/C _4524_/X vssd1 vssd1 vccd1 vccd1 _4526_/B sky130_fd_sc_hd__o21ai_1
X_8293_ _8359_/A _8359_/B _8291_/A vssd1 vssd1 vccd1 vccd1 _8293_/Y sky130_fd_sc_hd__o21ai_1
X_4456_ _5049_/A vssd1 vssd1 vccd1 vccd1 _5132_/A sky130_fd_sc_hd__clkbuf_2
X_7244_ _7244_/A _7244_/B vssd1 vssd1 vccd1 vccd1 _7253_/B sky130_fd_sc_hd__nor2_1
X_4387_ _4387_/A vssd1 vssd1 vccd1 vccd1 _4387_/Y sky130_fd_sc_hd__clkinv_2
X_7175_ _7180_/A _7175_/B vssd1 vssd1 vccd1 vccd1 _7206_/B sky130_fd_sc_hd__nor2_1
X_6126_ _6126_/A _6126_/B vssd1 vssd1 vccd1 vccd1 _6184_/B sky130_fd_sc_hd__and2_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6057_ _6057_/A _6057_/B vssd1 vssd1 vccd1 vccd1 _6059_/B sky130_fd_sc_hd__xor2_1
XFILLER_45_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5008_ _5035_/D _5092_/B _4996_/B _4972_/A _5012_/A vssd1 vssd1 vccd1 vccd1 _5009_/D
+ sky130_fd_sc_hd__o41a_1
XFILLER_26_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6959_ _6910_/B _6955_/Y _6954_/A _6954_/Y vssd1 vssd1 vccd1 vccd1 _6960_/C sky130_fd_sc_hd__a211o_1
XFILLER_5_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4310_ _4314_/A vssd1 vssd1 vccd1 vccd1 _4310_/Y sky130_fd_sc_hd__inv_2
X_5290_ _8504_/Q _5290_/B vssd1 vssd1 vccd1 vccd1 _5291_/C sky130_fd_sc_hd__nand2_1
XFILLER_67_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7931_ _7993_/A _7931_/B vssd1 vssd1 vccd1 vccd1 _7934_/A sky130_fd_sc_hd__nand2_1
XFILLER_63_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7862_ _7945_/A _7862_/B vssd1 vssd1 vccd1 vccd1 _7864_/C sky130_fd_sc_hd__xnor2_1
XFILLER_23_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6813_ _6839_/A _6812_/C _6812_/A vssd1 vssd1 vccd1 vccd1 _6814_/C sky130_fd_sc_hd__a21o_1
X_7793_ _7792_/B _7792_/C _7792_/A vssd1 vssd1 vccd1 vccd1 _7795_/B sky130_fd_sc_hd__o21ai_1
X_6744_ _6914_/B vssd1 vssd1 vccd1 vccd1 _6980_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_23_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6675_ _6675_/A _6698_/A vssd1 vssd1 vccd1 vccd1 _6703_/A sky130_fd_sc_hd__nand2_1
X_5626_ _5628_/A _5627_/A vssd1 vssd1 vccd1 vccd1 _5754_/A sky130_fd_sc_hd__or2_2
X_8414_ _8406_/B _8414_/B vssd1 vssd1 vccd1 vccd1 _8415_/C sky130_fd_sc_hd__and2b_1
X_8345_ _8345_/A _8288_/A vssd1 vssd1 vccd1 vccd1 _8345_/X sky130_fd_sc_hd__or2b_1
X_5557_ _5557_/A _5677_/A _5557_/C vssd1 vssd1 vccd1 vccd1 _5677_/B sky130_fd_sc_hd__nor3_1
X_4508_ _8453_/Q _5325_/B vssd1 vssd1 vccd1 vccd1 _5327_/B sky130_fd_sc_hd__nand2_1
X_8276_ _8277_/A _8276_/B _8276_/C vssd1 vssd1 vccd1 vccd1 _8278_/A sky130_fd_sc_hd__and3b_1
XFILLER_2_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5488_ _5488_/A vssd1 vssd1 vccd1 vccd1 _5488_/Y sky130_fd_sc_hd__inv_2
X_7227_ _7226_/A _7226_/C _7226_/B vssd1 vssd1 vccd1 vccd1 _7228_/C sky130_fd_sc_hd__o21a_1
X_4439_ _8473_/Q vssd1 vssd1 vccd1 vccd1 _7644_/B sky130_fd_sc_hd__inv_2
X_7158_ _7193_/A _7193_/B vssd1 vssd1 vccd1 vccd1 _7173_/B sky130_fd_sc_hd__xor2_1
XFILLER_76_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7089_ _7021_/Y _7022_/X _7017_/B _7019_/C vssd1 vssd1 vccd1 vccd1 _7089_/Y sky130_fd_sc_hd__o211ai_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6109_ _6110_/A _6110_/B _6110_/C vssd1 vssd1 vccd1 vccd1 _6111_/A sky130_fd_sc_hd__o21a_1
XFILLER_27_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8622__38 vssd1 vssd1 vccd1 vccd1 _8622__38/HI _8717_/A sky130_fd_sc_hd__conb_1
XFILLER_18_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4790_ _4790_/A _4790_/B _4953_/B vssd1 vssd1 vccd1 vccd1 _5055_/A sky130_fd_sc_hd__nor3_4
XFILLER_20_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6460_ _6459_/A _6466_/A _6466_/B _6459_/D vssd1 vssd1 vccd1 vccd1 _6461_/B sky130_fd_sc_hd__a22oi_1
X_6391_ _8567_/Q vssd1 vssd1 vccd1 vccd1 _7410_/A sky130_fd_sc_hd__clkinv_2
X_5411_ _5705_/A _5410_/A _5860_/A _5410_/Y vssd1 vssd1 vccd1 vccd1 _5412_/B sky130_fd_sc_hd__o31a_1
X_8130_ _8131_/A _8131_/B vssd1 vssd1 vccd1 vccd1 _8132_/A sky130_fd_sc_hd__nand2_1
X_5342_ _5374_/A _5337_/B _5336_/A vssd1 vssd1 vccd1 vccd1 _5343_/B sky130_fd_sc_hd__o21a_1
X_8061_ _8260_/C _7844_/Y _7964_/A _7964_/B vssd1 vssd1 vccd1 vccd1 _8066_/A sky130_fd_sc_hd__a22o_1
X_7012_ _6947_/A _7079_/B _7011_/Y vssd1 vssd1 vccd1 vccd1 _7017_/A sky130_fd_sc_hd__o21ai_2
X_5273_ _5273_/A vssd1 vssd1 vccd1 vccd1 _8498_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7914_ _7914_/A _8231_/A vssd1 vssd1 vccd1 vccd1 _8299_/A sky130_fd_sc_hd__xor2_4
XFILLER_63_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7845_ _7742_/A _7885_/B _7885_/C _7844_/A _7725_/C vssd1 vssd1 vccd1 vccd1 _7845_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_36_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4988_ _5092_/A _4939_/B _4987_/X _4839_/A vssd1 vssd1 vccd1 vccd1 _4988_/X sky130_fd_sc_hd__o31a_1
X_7776_ _7660_/A _7660_/B _7546_/A _7526_/B vssd1 vssd1 vccd1 vccd1 _7778_/B sky130_fd_sc_hd__o2bb2a_1
X_6727_ _6727_/A _6727_/B vssd1 vssd1 vccd1 vccd1 _6729_/B sky130_fd_sc_hd__xnor2_1
X_6658_ _6658_/A _6678_/B vssd1 vssd1 vccd1 vccd1 _6660_/B sky130_fd_sc_hd__xnor2_1
X_5609_ _5609_/A _5609_/B _5609_/C vssd1 vssd1 vccd1 vccd1 _5722_/A sky130_fd_sc_hd__or3_1
X_6589_ _8555_/Q vssd1 vssd1 vccd1 vccd1 _6590_/A sky130_fd_sc_hd__inv_2
XFILLER_11_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8328_ _8069_/A _8274_/S _8273_/Y vssd1 vssd1 vccd1 vccd1 _8329_/B sky130_fd_sc_hd__o21a_1
XFILLER_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8259_ _8152_/A _8152_/B _8258_/X vssd1 vssd1 vccd1 vccd1 _8266_/A sky130_fd_sc_hd__o21ai_1
XFILLER_78_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5960_ _5963_/A _5963_/B vssd1 vssd1 vccd1 vccd1 _5961_/B sky130_fd_sc_hd__xor2_1
X_4911_ _5049_/A _5151_/C _4955_/B _5020_/C vssd1 vssd1 vccd1 vccd1 _4911_/X sky130_fd_sc_hd__or4_1
XFILLER_80_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5891_ _5893_/A _5893_/B vssd1 vssd1 vccd1 vccd1 _6067_/A sky130_fd_sc_hd__and2_1
X_7630_ _8147_/A vssd1 vssd1 vccd1 vccd1 _8326_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_33_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4842_ _5031_/B _4993_/A _4842_/C vssd1 vssd1 vccd1 vccd1 _4842_/X sky130_fd_sc_hd__or3_1
XFILLER_20_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4773_ _4773_/A vssd1 vssd1 vccd1 vccd1 _4786_/B sky130_fd_sc_hd__clkbuf_2
X_7561_ _8405_/A _7553_/B _7574_/A _7574_/B _7556_/A vssd1 vssd1 vccd1 vccd1 _7562_/C
+ sky130_fd_sc_hd__a221o_1
X_6512_ _6512_/A _6512_/B vssd1 vssd1 vccd1 vccd1 _6570_/A sky130_fd_sc_hd__nor2_1
X_7492_ _8467_/Q _8570_/Q vssd1 vssd1 vccd1 vccd1 _7493_/A sky130_fd_sc_hd__or2b_1
X_6443_ _6439_/A _5294_/X _6432_/X _6442_/X vssd1 vssd1 vccd1 vccd1 _8552_/D sky130_fd_sc_hd__a22o_1
X_6374_ _6374_/A vssd1 vssd1 vccd1 vccd1 _8541_/D sky130_fd_sc_hd__clkbuf_1
X_5325_ _8453_/Q _5325_/B vssd1 vssd1 vccd1 vccd1 _5326_/B sky130_fd_sc_hd__and2_2
X_8113_ _8113_/A _8113_/B vssd1 vssd1 vccd1 vccd1 _8114_/B sky130_fd_sc_hd__xnor2_2
X_5256_ _6396_/D _5258_/C _5230_/B vssd1 vssd1 vccd1 vccd1 _5256_/Y sky130_fd_sc_hd__o21ai_1
X_8044_ _8127_/A _8044_/B vssd1 vssd1 vccd1 vccd1 _8045_/B sky130_fd_sc_hd__and2_1
XFILLER_87_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5187_ _5131_/X _5186_/X _5207_/A vssd1 vssd1 vccd1 vccd1 _5202_/A sky130_fd_sc_hd__o21ai_2
XFILLER_68_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7828_ _7978_/A vssd1 vssd1 vccd1 vccd1 _7984_/A sky130_fd_sc_hd__clkinv_2
X_7759_ _7837_/B _7758_/C _7758_/A vssd1 vssd1 vccd1 vccd1 _7788_/B sky130_fd_sc_hd__a21o_1
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5110_ _5110_/A _5118_/B vssd1 vssd1 vccd1 vccd1 _5110_/X sky130_fd_sc_hd__or2_1
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6090_ _6087_/A _6090_/B _6090_/C _6090_/D vssd1 vssd1 vccd1 vccd1 _6090_/X sky130_fd_sc_hd__and4b_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5041_ _5162_/A _5148_/A _5041_/C _5071_/C vssd1 vssd1 vccd1 vccd1 _5041_/X sky130_fd_sc_hd__or4_1
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8731_ _8731_/A _4317_/Y vssd1 vssd1 vccd1 vccd1 io_out[16] sky130_fd_sc_hd__ebufn_8
XFILLER_80_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6992_ _6992_/A _6992_/B vssd1 vssd1 vccd1 vccd1 _6993_/B sky130_fd_sc_hd__xor2_1
XFILLER_53_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5943_ _5943_/A _5943_/B vssd1 vssd1 vccd1 vccd1 _6015_/B sky130_fd_sc_hd__xor2_1
X_5874_ _5812_/A _5812_/B _5813_/A vssd1 vssd1 vccd1 vccd1 _5887_/A sky130_fd_sc_hd__a21oi_1
XFILLER_33_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4825_ _5064_/B _5064_/D vssd1 vssd1 vccd1 vccd1 _5051_/A sky130_fd_sc_hd__or2_2
X_7613_ _7416_/X _7613_/B vssd1 vssd1 vccd1 vccd1 _7613_/X sky130_fd_sc_hd__and2b_1
XFILLER_21_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7544_ _8367_/A _7803_/A vssd1 vssd1 vccd1 vccd1 _7639_/A sky130_fd_sc_hd__nand2_1
X_4756_ _4756_/A vssd1 vssd1 vccd1 vccd1 _4908_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_4687_ _5380_/B vssd1 vssd1 vccd1 vccd1 _7501_/B sky130_fd_sc_hd__inv_2
X_7475_ _7507_/A _7482_/B _7474_/X vssd1 vssd1 vccd1 vccd1 _7477_/C sky130_fd_sc_hd__a21oi_1
X_6426_ _6426_/A _6426_/B vssd1 vssd1 vccd1 vccd1 _8549_/D sky130_fd_sc_hd__nand2_1
X_6357_ _8536_/Q _8535_/Q _6357_/C vssd1 vssd1 vccd1 vccd1 _6362_/C sky130_fd_sc_hd__and3_1
X_8658__74 vssd1 vssd1 vccd1 vccd1 _8658__74/HI _8767_/A sky130_fd_sc_hd__conb_1
X_5308_ _6281_/B vssd1 vssd1 vccd1 vccd1 _6293_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6288_ _6289_/A _6289_/B _6289_/C _6289_/D vssd1 vssd1 vccd1 vccd1 _6288_/Y sky130_fd_sc_hd__o22ai_1
XFILLER_0_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5239_ _5239_/A vssd1 vssd1 vccd1 vccd1 _8488_/D sky130_fd_sc_hd__clkbuf_1
X_8027_ _8299_/A _8093_/B vssd1 vssd1 vccd1 vccd1 _8028_/B sky130_fd_sc_hd__xor2_1
XFILLER_29_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4610_ _4619_/A _4619_/B vssd1 vssd1 vccd1 vccd1 _4612_/B sky130_fd_sc_hd__nand2_1
XFILLER_30_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5590_ _5590_/A vssd1 vssd1 vccd1 vccd1 _6082_/B sky130_fd_sc_hd__inv_2
X_4541_ _4543_/B _4568_/B _4541_/C vssd1 vssd1 vccd1 vccd1 _4542_/A sky130_fd_sc_hd__and3b_1
X_7260_ _7217_/Y _7344_/B _7258_/Y _7343_/A vssd1 vssd1 vccd1 vccd1 _7338_/C sky130_fd_sc_hd__a211o_1
X_4472_ _8474_/Q _4480_/B vssd1 vssd1 vccd1 vccd1 _4473_/A sky130_fd_sc_hd__and2_1
X_7191_ _7191_/A _7191_/B vssd1 vssd1 vccd1 vccd1 _7212_/B sky130_fd_sc_hd__xnor2_1
X_6211_ _6211_/A _6211_/B vssd1 vssd1 vccd1 vccd1 _6211_/Y sky130_fd_sc_hd__nand2_1
X_6142_ _6143_/A _6143_/B vssd1 vssd1 vccd1 vccd1 _6144_/A sky130_fd_sc_hd__nand2_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6073_ _6073_/A _6073_/B vssd1 vssd1 vccd1 vccd1 _6073_/X sky130_fd_sc_hd__or2_1
X_5024_ _5121_/A vssd1 vssd1 vccd1 vccd1 _5080_/A sky130_fd_sc_hd__clkbuf_2
XINSDIODE2_29 _8710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_18 _8705_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6975_ _7034_/S _6975_/B vssd1 vssd1 vccd1 vccd1 _6975_/X sky130_fd_sc_hd__and2_1
XFILLER_65_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8714_ _8714_/A _4297_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[31] sky130_fd_sc_hd__ebufn_8
X_5926_ _5853_/A _5853_/B _5925_/X vssd1 vssd1 vccd1 vccd1 _5956_/A sky130_fd_sc_hd__a21oi_2
XFILLER_34_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5857_ _5861_/A _5800_/B _5861_/C vssd1 vssd1 vccd1 vccd1 _5857_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_21_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4808_ _4808_/A _4809_/B vssd1 vssd1 vccd1 vccd1 _5112_/A sky130_fd_sc_hd__nor2_2
XFILLER_21_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5788_ _5788_/A _5788_/B vssd1 vssd1 vccd1 vccd1 _5818_/B sky130_fd_sc_hd__xor2_2
X_8576_ input3/X _8576_/D vssd1 vssd1 vccd1 vccd1 _8576_/Q sky130_fd_sc_hd__dfxtp_1
X_4739_ _5144_/C _5144_/B vssd1 vssd1 vccd1 vccd1 _4742_/B sky130_fd_sc_hd__xnor2_1
X_7527_ _7813_/A _7695_/B _7528_/C vssd1 vssd1 vccd1 vccd1 _7655_/A sky130_fd_sc_hd__a21oi_1
XFILLER_79_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7458_ _8569_/Q _7501_/A vssd1 vssd1 vccd1 vccd1 _7459_/B sky130_fd_sc_hd__and2b_1
X_6409_ _8567_/Q _6424_/B _6409_/C vssd1 vssd1 vccd1 vccd1 _6409_/X sky130_fd_sc_hd__or3_1
X_7389_ _7384_/B _5241_/X _6432_/X _7388_/X vssd1 vssd1 vccd1 vccd1 _8563_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6760_ _6558_/A _6721_/A _6679_/B vssd1 vssd1 vccd1 vccd1 _7026_/A sky130_fd_sc_hd__o21ai_4
XFILLER_50_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5711_ _5805_/A _5711_/B vssd1 vssd1 vccd1 vccd1 _5711_/Y sky130_fd_sc_hd__nor2_1
X_6691_ _6791_/A _6691_/B vssd1 vssd1 vccd1 vccd1 _6777_/B sky130_fd_sc_hd__nor2_1
X_5642_ _5684_/A _5650_/A vssd1 vssd1 vccd1 vccd1 _5976_/A sky130_fd_sc_hd__nand2_1
X_8430_ _8430_/A _8430_/B vssd1 vssd1 vccd1 vccd1 _8430_/Y sky130_fd_sc_hd__nor2_1
XFILLER_31_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5573_ _5574_/A _5574_/B vssd1 vssd1 vccd1 vccd1 _5575_/A sky130_fd_sc_hd__nor2_1
X_8361_ _8361_/A _8361_/B vssd1 vssd1 vccd1 vccd1 _8362_/C sky130_fd_sc_hd__xnor2_1
X_7312_ _7312_/A _7312_/B vssd1 vssd1 vccd1 vccd1 _7313_/B sky130_fd_sc_hd__xnor2_1
X_4524_ _4568_/B vssd1 vssd1 vccd1 vccd1 _4524_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_8292_ _8292_/A vssd1 vssd1 vccd1 vccd1 _8359_/A sky130_fd_sc_hd__inv_2
X_4455_ _5064_/A _4945_/A vssd1 vssd1 vccd1 vccd1 _5049_/A sky130_fd_sc_hd__or2_1
X_7243_ _7243_/A _7243_/B vssd1 vssd1 vccd1 vccd1 _7349_/A sky130_fd_sc_hd__nor2_1
X_7174_ _7155_/A _7155_/C _7155_/B vssd1 vssd1 vccd1 vccd1 _7177_/B sky130_fd_sc_hd__a21o_1
X_4386_ _4387_/A vssd1 vssd1 vccd1 vccd1 _4386_/Y sky130_fd_sc_hd__inv_2
X_8628__44 vssd1 vssd1 vccd1 vccd1 _8628__44/HI _8723_/A sky130_fd_sc_hd__conb_1
XFILLER_58_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6125_ _6125_/A _6125_/B vssd1 vssd1 vccd1 vccd1 _6132_/B sky130_fd_sc_hd__and2_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6056_ _5669_/B _5669_/C _5669_/A vssd1 vssd1 vccd1 vccd1 _6058_/A sky130_fd_sc_hd__a21boi_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5007_ _5064_/B _5012_/C vssd1 vssd1 vccd1 vccd1 _5092_/B sky130_fd_sc_hd__or2_1
XFILLER_66_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6958_ _6953_/A _6953_/B _6957_/X vssd1 vssd1 vccd1 vccd1 _6960_/B sky130_fd_sc_hd__a21o_1
XFILLER_81_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6889_ _6888_/A _6889_/B vssd1 vssd1 vccd1 vccd1 _7277_/A sky130_fd_sc_hd__and2b_1
X_5909_ _5708_/X _5882_/B _5880_/Y vssd1 vssd1 vccd1 vccd1 _5911_/B sky130_fd_sc_hd__a21oi_2
XFILLER_22_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8559_ input3/X _8559_/D vssd1 vssd1 vccd1 vccd1 _8559_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7930_ _7930_/A _7930_/B _7930_/C vssd1 vssd1 vccd1 vccd1 _7931_/B sky130_fd_sc_hd__nand3_1
XFILLER_82_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7861_ _7861_/A _7886_/A vssd1 vssd1 vccd1 vccd1 _7862_/B sky130_fd_sc_hd__xnor2_1
X_6812_ _6812_/A _6839_/A _6812_/C vssd1 vssd1 vccd1 vccd1 _6839_/B sky130_fd_sc_hd__nand3_1
XFILLER_35_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7792_ _7792_/A _7792_/B _7792_/C vssd1 vssd1 vccd1 vccd1 _8193_/B sky130_fd_sc_hd__or3_1
X_6743_ _6816_/A _6742_/C _6829_/A vssd1 vssd1 vccd1 vccd1 _6758_/C sky130_fd_sc_hd__a21o_1
X_6674_ _6780_/A _6675_/A _6674_/C vssd1 vssd1 vccd1 vccd1 _6698_/A sky130_fd_sc_hd__nand3_1
X_5625_ _5625_/A _5625_/B vssd1 vssd1 vccd1 vccd1 _5631_/B sky130_fd_sc_hd__nand2_1
X_8413_ _8421_/A _8413_/B vssd1 vssd1 vccd1 vccd1 _8415_/B sky130_fd_sc_hd__or2_1
X_8344_ _8344_/A _8344_/B vssd1 vssd1 vccd1 vccd1 _8351_/A sky130_fd_sc_hd__xnor2_2
X_5556_ _5555_/B _5555_/C _5561_/A vssd1 vssd1 vccd1 vccd1 _5557_/C sky130_fd_sc_hd__a21oi_1
X_8275_ _8326_/C _8275_/B vssd1 vssd1 vccd1 vccd1 _8279_/A sky130_fd_sc_hd__xor2_2
X_5487_ _5492_/B _5488_/A vssd1 vssd1 vccd1 vccd1 _5487_/X sky130_fd_sc_hd__xor2_2
X_4507_ _8441_/Q _4507_/B _4507_/C vssd1 vssd1 vccd1 vccd1 _5325_/B sky130_fd_sc_hd__or3_1
X_7226_ _7226_/A _7226_/B _7226_/C vssd1 vssd1 vccd1 vccd1 _7228_/B sky130_fd_sc_hd__nor3_1
X_4438_ _4438_/A _4467_/C vssd1 vssd1 vccd1 vccd1 _4438_/Y sky130_fd_sc_hd__nor2_1
X_7157_ _7177_/A _7159_/B vssd1 vssd1 vccd1 vccd1 _7173_/A sky130_fd_sc_hd__xnor2_1
X_4369_ _4369_/A vssd1 vssd1 vccd1 vccd1 _4369_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7088_ _7143_/A _7143_/B _7143_/C vssd1 vssd1 vccd1 vccd1 _7088_/Y sky130_fd_sc_hd__nor3_1
XFILLER_58_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6108_ _6108_/A _6108_/B vssd1 vssd1 vccd1 vccd1 _6110_/C sky130_fd_sc_hd__xor2_1
XFILLER_86_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6039_ _6160_/A _6160_/B vssd1 vssd1 vccd1 vccd1 _6040_/B sky130_fd_sc_hd__xor2_1
XFILLER_26_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6390_ _6390_/A vssd1 vssd1 vccd1 vccd1 _8547_/D sky130_fd_sc_hd__clkbuf_1
X_5410_ _5410_/A _5565_/A vssd1 vssd1 vccd1 vccd1 _5410_/Y sky130_fd_sc_hd__nand2_1
X_5341_ _5341_/A _5341_/B vssd1 vssd1 vccd1 vccd1 _5343_/A sky130_fd_sc_hd__nor2_1
X_8060_ _8317_/A _8147_/B vssd1 vssd1 vccd1 vccd1 _8260_/C sky130_fd_sc_hd__nor2_2
X_5272_ _5277_/C _5291_/A _5272_/C vssd1 vssd1 vccd1 vccd1 _5273_/A sky130_fd_sc_hd__and3b_1
X_7011_ _7075_/A _7011_/B vssd1 vssd1 vccd1 vccd1 _7011_/Y sky130_fd_sc_hd__nand2_1
XFILLER_68_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7913_ _7913_/A vssd1 vssd1 vccd1 vccd1 _8231_/A sky130_fd_sc_hd__buf_2
XFILLER_51_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7844_ _7844_/A _8146_/A _8146_/B vssd1 vssd1 vccd1 vccd1 _7844_/Y sky130_fd_sc_hd__nor3_2
XFILLER_24_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7775_ _7818_/A _7818_/B vssd1 vssd1 vccd1 vccd1 _7781_/A sky130_fd_sc_hd__xnor2_1
X_4987_ _4987_/A _5117_/B vssd1 vssd1 vccd1 vccd1 _4987_/X sky130_fd_sc_hd__or2_1
X_6726_ _6937_/B _6937_/C _6937_/A vssd1 vssd1 vccd1 vccd1 _6729_/A sky130_fd_sc_hd__a21boi_1
XFILLER_51_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6657_ _6657_/A _6657_/B vssd1 vssd1 vccd1 vccd1 _6678_/B sky130_fd_sc_hd__xnor2_4
X_6588_ _6543_/X _6604_/A _6596_/B _6595_/A vssd1 vssd1 vccd1 vccd1 _6592_/A sky130_fd_sc_hd__a31o_1
X_5608_ _5615_/A _5488_/A _5609_/C _5764_/A vssd1 vssd1 vccd1 vccd1 _5610_/B sky130_fd_sc_hd__o22ai_1
XFILLER_3_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5539_ _5539_/A _5539_/B vssd1 vssd1 vccd1 vccd1 _5547_/A sky130_fd_sc_hd__xnor2_1
X_8327_ _7618_/A _7618_/C _7615_/B vssd1 vssd1 vccd1 vccd1 _8329_/A sky130_fd_sc_hd__a21oi_1
XFILLER_11_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8258_ _8258_/A _8258_/B vssd1 vssd1 vccd1 vccd1 _8258_/X sky130_fd_sc_hd__or2_1
XFILLER_78_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7209_ _7219_/A _7219_/B _7206_/X _7180_/C vssd1 vssd1 vccd1 vccd1 _7211_/B sky130_fd_sc_hd__o2bb2a_1
X_8189_ _8201_/A _8201_/B _8201_/C vssd1 vssd1 vccd1 vccd1 _8202_/A sky130_fd_sc_hd__o21a_1
XFILLER_54_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4910_ _4910_/A vssd1 vssd1 vccd1 vccd1 _5020_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_92_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5890_ _5890_/A _5890_/B vssd1 vssd1 vccd1 vccd1 _5893_/B sky130_fd_sc_hd__xor2_1
XFILLER_18_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4841_ _4960_/A _5011_/A vssd1 vssd1 vccd1 vccd1 _4842_/C sky130_fd_sc_hd__or2_1
XFILLER_60_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4772_ _4772_/A _4909_/B _4771_/X vssd1 vssd1 vccd1 vccd1 _4897_/A sky130_fd_sc_hd__or3b_1
XFILLER_20_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7560_ _7569_/A _7569_/B _7559_/X vssd1 vssd1 vccd1 vccd1 _7574_/B sky130_fd_sc_hd__a21o_2
X_6511_ _7410_/A _7613_/B vssd1 vssd1 vccd1 vccd1 _6512_/B sky130_fd_sc_hd__nor2_1
XFILLER_9_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7491_ _7766_/A _7489_/Y _7490_/Y vssd1 vssd1 vccd1 vccd1 _8576_/D sky130_fd_sc_hd__a21oi_1
X_6442_ _6442_/A _6442_/B vssd1 vssd1 vccd1 vccd1 _6442_/X sky130_fd_sc_hd__xor2_1
X_6373_ _6375_/B _6389_/B _6373_/C vssd1 vssd1 vccd1 vccd1 _6374_/A sky130_fd_sc_hd__and3b_1
X_8112_ _8110_/Y _8112_/B vssd1 vssd1 vccd1 vccd1 _8113_/B sky130_fd_sc_hd__and2b_1
X_5324_ _5322_/C _5318_/Y _5323_/X _5213_/X vssd1 vssd1 vccd1 vccd1 _8508_/D sky130_fd_sc_hd__o211a_1
X_5255_ _5258_/C _5255_/B vssd1 vssd1 vccd1 vccd1 _8493_/D sky130_fd_sc_hd__nor2_1
X_8043_ _8127_/A _8044_/B vssd1 vssd1 vccd1 vccd1 _8131_/A sky130_fd_sc_hd__nor2_1
X_5186_ _4711_/A _5178_/B _5046_/Y _5176_/X _5185_/Y vssd1 vssd1 vccd1 vccd1 _5186_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_28_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7827_ _8367_/B _7808_/A _7825_/A vssd1 vssd1 vccd1 vccd1 _7827_/X sky130_fd_sc_hd__a21o_1
XFILLER_12_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7758_ _7758_/A _7837_/B _7758_/C vssd1 vssd1 vccd1 vccd1 _7788_/A sky130_fd_sc_hd__nand3_1
X_6709_ _6731_/A _6731_/B vssd1 vssd1 vccd1 vccd1 _6907_/A sky130_fd_sc_hd__xnor2_1
X_7689_ _7690_/A _7690_/B vssd1 vssd1 vccd1 vccd1 _7691_/A sky130_fd_sc_hd__nor2_1
XFILLER_3_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5040_ _5148_/B _5040_/B _5169_/B vssd1 vssd1 vccd1 vccd1 _5118_/A sky130_fd_sc_hd__or3_1
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6991_ _6991_/A _6991_/B vssd1 vssd1 vccd1 vccd1 _6992_/B sky130_fd_sc_hd__and2_1
XFILLER_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8730_ _8730_/A _4316_/Y vssd1 vssd1 vccd1 vccd1 io_out[15] sky130_fd_sc_hd__ebufn_8
XFILLER_65_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5942_ _5949_/A _5942_/B vssd1 vssd1 vccd1 vccd1 _5943_/B sky130_fd_sc_hd__xnor2_1
XFILLER_80_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5873_ _5873_/A _5896_/B vssd1 vssd1 vccd1 vccd1 _5890_/A sky130_fd_sc_hd__xnor2_1
X_4824_ _4960_/A _4968_/A _5171_/C _5090_/B vssd1 vssd1 vccd1 vccd1 _5064_/D sky130_fd_sc_hd__nor4_1
X_7612_ _7612_/A vssd1 vssd1 vccd1 vccd1 _7618_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4755_ _4755_/A _4765_/A _5144_/C vssd1 vssd1 vccd1 vccd1 _4756_/A sky130_fd_sc_hd__nor3b_1
XFILLER_21_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7543_ _7649_/A _7649_/B vssd1 vssd1 vccd1 vccd1 _7803_/A sky130_fd_sc_hd__xor2_4
X_4686_ _4686_/A vssd1 vssd1 vccd1 vccd1 _8468_/D sky130_fd_sc_hd__clkbuf_1
X_7474_ _7507_/A _7482_/B _7467_/X vssd1 vssd1 vccd1 vccd1 _7474_/X sky130_fd_sc_hd__o21a_1
X_6425_ _6424_/B _6422_/Y _6424_/X _6450_/B vssd1 vssd1 vccd1 vccd1 _6426_/B sky130_fd_sc_hd__a2bb2o_1
X_6356_ _6356_/A _6356_/B vssd1 vssd1 vccd1 vccd1 _8535_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5307_ _8526_/Q vssd1 vssd1 vccd1 vccd1 _5495_/A sky130_fd_sc_hd__inv_2
X_8673__89 vssd1 vssd1 vccd1 vccd1 _8673__89/HI _8782_/A sky130_fd_sc_hd__conb_1
X_8026_ _8231_/A _7980_/Y _8025_/X vssd1 vssd1 vccd1 vccd1 _8093_/B sky130_fd_sc_hd__o21a_1
X_6287_ _6286_/B _6293_/B vssd1 vssd1 vccd1 vccd1 _6289_/D sky130_fd_sc_hd__and2b_1
X_5238_ _5240_/B _5291_/A _5238_/C vssd1 vssd1 vccd1 vccd1 _5239_/A sky130_fd_sc_hd__and3b_1
XFILLER_75_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5169_ _5169_/A _5169_/B _5169_/C _5169_/D vssd1 vssd1 vccd1 vccd1 _5169_/X sky130_fd_sc_hd__or4_1
XFILLER_29_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4540_ _8440_/Q _4539_/C _8441_/Q vssd1 vssd1 vccd1 vccd1 _4541_/C sky130_fd_sc_hd__a21o_1
X_4471_ _4495_/B vssd1 vssd1 vccd1 vccd1 _4480_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_7_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7190_ _7185_/A _7185_/B _7186_/A _7182_/B _7205_/A vssd1 vssd1 vccd1 vccd1 _7212_/A
+ sky130_fd_sc_hd__o32ai_4
X_6210_ _6210_/A _6210_/B vssd1 vssd1 vccd1 vccd1 _6213_/A sky130_fd_sc_hd__xnor2_1
X_6141_ _6141_/A _6141_/B vssd1 vssd1 vccd1 vccd1 _6143_/B sky130_fd_sc_hd__xnor2_1
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6072_ _6073_/A _6073_/B vssd1 vssd1 vccd1 vccd1 _6084_/B sky130_fd_sc_hd__xnor2_1
XINSDIODE2_19 _8705_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5023_ _4619_/A _5017_/X _5022_/X _5175_/S vssd1 vssd1 vccd1 vccd1 _5023_/X sky130_fd_sc_hd__o211a_1
XFILLER_57_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6974_ _6745_/B _7044_/A _7044_/B _7176_/B vssd1 vssd1 vccd1 vccd1 _6975_/B sky130_fd_sc_hd__a31o_1
XFILLER_26_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8713_ _8713_/A _4295_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[30] sky130_fd_sc_hd__ebufn_8
X_5925_ _5925_/A _5925_/B vssd1 vssd1 vccd1 vccd1 _5925_/X sky130_fd_sc_hd__and2_1
XFILLER_41_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5856_ _5901_/A vssd1 vssd1 vccd1 vccd1 _5999_/A sky130_fd_sc_hd__inv_2
XFILLER_21_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4807_ _4993_/B _4993_/A vssd1 vssd1 vccd1 vccd1 _4969_/B sky130_fd_sc_hd__or2_1
X_5787_ _5932_/B _5785_/Y _5868_/A vssd1 vssd1 vccd1 vccd1 _5788_/B sky130_fd_sc_hd__a21oi_2
X_8575_ input3/X _8575_/D vssd1 vssd1 vccd1 vccd1 _8575_/Q sky130_fd_sc_hd__dfxtp_1
X_4738_ _5380_/B _4738_/B vssd1 vssd1 vccd1 vccd1 _5144_/B sky130_fd_sc_hd__nor2_1
X_7526_ _7770_/A _7526_/B vssd1 vssd1 vccd1 vccd1 _7528_/C sky130_fd_sc_hd__nor2_1
X_4669_ _4735_/B _4661_/B _5192_/B _4790_/A _4668_/X vssd1 vssd1 vccd1 vccd1 _8465_/D
+ sky130_fd_sc_hd__o221a_1
X_7457_ _7457_/A vssd1 vssd1 vccd1 vccd1 _8571_/D sky130_fd_sc_hd__clkbuf_1
X_6408_ _7384_/B _7380_/A _6562_/B vssd1 vssd1 vccd1 vccd1 _6409_/C sky130_fd_sc_hd__o21a_1
X_7388_ _7388_/A _7388_/B vssd1 vssd1 vccd1 vccd1 _7388_/X sky130_fd_sc_hd__xor2_1
XFILLER_1_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6339_ _6343_/C _6339_/B _6382_/B vssd1 vssd1 vccd1 vccd1 _6340_/A sky130_fd_sc_hd__and3b_1
XFILLER_0_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8009_ _8010_/A _8010_/B vssd1 vssd1 vccd1 vccd1 _8011_/A sky130_fd_sc_hd__nand2_1
XFILLER_29_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5710_ _5805_/A _5711_/B _5707_/Y _5708_/X _5861_/A vssd1 vssd1 vccd1 vccd1 _5914_/A
+ sky130_fd_sc_hd__o2111a_1
X_6690_ _6690_/A _7294_/B _6690_/C vssd1 vssd1 vccd1 vccd1 _6691_/B sky130_fd_sc_hd__nor3_1
XFILLER_31_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5641_ _5664_/A _5664_/B vssd1 vssd1 vccd1 vccd1 _5699_/A sky130_fd_sc_hd__or2_1
X_8360_ _8359_/A _8359_/B _8359_/C vssd1 vssd1 vccd1 vccd1 _8362_/B sky130_fd_sc_hd__a21o_1
X_5572_ _5466_/A _5831_/A _5586_/A _5586_/B vssd1 vssd1 vccd1 vccd1 _5574_/B sky130_fd_sc_hd__o22a_1
X_7311_ _6828_/A _6828_/B _6825_/Y vssd1 vssd1 vccd1 vccd1 _7312_/B sky130_fd_sc_hd__a21oi_1
X_4523_ _4536_/A vssd1 vssd1 vccd1 vccd1 _4568_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_8291_ _8291_/A _8291_/B vssd1 vssd1 vccd1 vccd1 _8359_/C sky130_fd_sc_hd__xnor2_1
X_7242_ _7241_/A _7241_/B _7241_/C vssd1 vssd1 vccd1 vccd1 _7243_/B sky130_fd_sc_hd__a21oi_1
X_4454_ _5099_/A vssd1 vssd1 vccd1 vccd1 _4945_/A sky130_fd_sc_hd__clkbuf_2
X_7173_ _7173_/A _7173_/B vssd1 vssd1 vccd1 vccd1 _7191_/B sky130_fd_sc_hd__xnor2_1
X_4385_ _4387_/A vssd1 vssd1 vccd1 vccd1 _4385_/Y sky130_fd_sc_hd__inv_2
X_6124_ _6124_/A _6124_/B vssd1 vssd1 vccd1 vccd1 _6132_/A sky130_fd_sc_hd__nor2_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6055_ _6075_/A _6075_/B vssd1 vssd1 vccd1 vccd1 _6071_/A sky130_fd_sc_hd__xor2_1
X_8643__59 vssd1 vssd1 vccd1 vccd1 _8643__59/HI _8752_/A sky130_fd_sc_hd__conb_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5006_ _5109_/A _5109_/B _5006_/C _5006_/D vssd1 vssd1 vccd1 vccd1 _5006_/X sky130_fd_sc_hd__or4_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6957_ _6952_/A _6957_/B vssd1 vssd1 vccd1 vccd1 _6957_/X sky130_fd_sc_hd__and2b_1
XFILLER_81_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6888_ _6888_/A _6888_/B _6888_/C vssd1 vssd1 vccd1 vccd1 _6889_/B sky130_fd_sc_hd__or3_1
X_5908_ _5971_/A _5908_/B vssd1 vssd1 vccd1 vccd1 _5911_/A sky130_fd_sc_hd__xnor2_2
XFILLER_14_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5839_ _5839_/A _6137_/B vssd1 vssd1 vccd1 vccd1 _5841_/A sky130_fd_sc_hd__nor2_1
X_8558_ input3/X _8558_/D vssd1 vssd1 vccd1 vccd1 _8558_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7509_ _7680_/A _7680_/B vssd1 vssd1 vccd1 vccd1 _7921_/A sky130_fd_sc_hd__xnor2_4
X_8489_ input3/X _8489_/D vssd1 vssd1 vccd1 vccd1 _8489_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7860_ _7860_/A _7860_/B vssd1 vssd1 vccd1 vccd1 _7864_/B sky130_fd_sc_hd__and2_1
X_6811_ _6836_/A _7296_/A _7296_/B vssd1 vssd1 vccd1 vccd1 _6812_/C sky130_fd_sc_hd__or3_1
XFILLER_23_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7791_ _7788_/X _7789_/Y _7638_/A _7672_/B vssd1 vssd1 vccd1 vccd1 _7792_/C sky130_fd_sc_hd__o211a_1
X_6742_ _6812_/A _6816_/A _6742_/C vssd1 vssd1 vccd1 vccd1 _6816_/B sky130_fd_sc_hd__nand3_1
X_6673_ _6939_/B _7323_/B _7069_/B _7068_/B vssd1 vssd1 vccd1 vccd1 _6674_/C sky130_fd_sc_hd__o31ai_2
XFILLER_31_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5624_ _5825_/A _5839_/A _5624_/C vssd1 vssd1 vccd1 vccd1 _5631_/A sky130_fd_sc_hd__or3_1
X_8412_ _8428_/A _8412_/B vssd1 vssd1 vccd1 vccd1 _8413_/B sky130_fd_sc_hd__and2b_1
X_8343_ _8343_/A _8343_/B vssd1 vssd1 vccd1 vccd1 _8344_/B sky130_fd_sc_hd__xnor2_1
X_5555_ _5561_/A _5555_/B _5555_/C vssd1 vssd1 vccd1 vccd1 _5677_/A sky130_fd_sc_hd__and3_1
X_8274_ _7899_/X _8273_/Y _8274_/S vssd1 vssd1 vccd1 vccd1 _8275_/B sky130_fd_sc_hd__mux2_1
X_5486_ _5767_/A _5609_/C vssd1 vssd1 vccd1 vccd1 _5625_/A sky130_fd_sc_hd__nor2_2
X_4506_ _4516_/A _4506_/B _4506_/C _4506_/D vssd1 vssd1 vccd1 vccd1 _4507_/C sky130_fd_sc_hd__or4_1
X_7225_ _7211_/A _7211_/C _7211_/B vssd1 vssd1 vccd1 vccd1 _7226_/C sky130_fd_sc_hd__o21a_1
X_4437_ _4780_/A _4671_/A vssd1 vssd1 vccd1 vccd1 _4467_/C sky130_fd_sc_hd__and2_1
X_7156_ _7156_/A _7156_/B vssd1 vssd1 vccd1 vccd1 _7159_/B sky130_fd_sc_hd__xor2_1
XFILLER_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4368_ _4369_/A vssd1 vssd1 vccd1 vccd1 _4368_/Y sky130_fd_sc_hd__inv_2
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6107_ _6184_/A _6183_/S vssd1 vssd1 vccd1 vccd1 _6110_/A sky130_fd_sc_hd__nor2_1
X_4299_ _4301_/A vssd1 vssd1 vccd1 vccd1 _4299_/Y sky130_fd_sc_hd__inv_2
X_7087_ _7019_/Y _7083_/X _7082_/X _7065_/A vssd1 vssd1 vccd1 vccd1 _7143_/C sky130_fd_sc_hd__a211oi_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6038_ _5953_/A _5953_/B _6037_/X vssd1 vssd1 vccd1 vccd1 _6160_/B sky130_fd_sc_hd__a21oi_1
XFILLER_92_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7989_ _7989_/A _8252_/A vssd1 vssd1 vccd1 vccd1 _7990_/B sky130_fd_sc_hd__or2_1
XFILLER_25_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5340_ _5339_/B _5360_/B vssd1 vssd1 vccd1 vccd1 _5341_/B sky130_fd_sc_hd__and2b_1
X_5271_ _6392_/C _8496_/Q _5263_/B _8498_/Q vssd1 vssd1 vccd1 vccd1 _5272_/C sky130_fd_sc_hd__a31o_1
XFILLER_87_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7010_ _7075_/A _7011_/B vssd1 vssd1 vccd1 vccd1 _7079_/B sky130_fd_sc_hd__xnor2_1
XFILLER_68_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8613__29 vssd1 vssd1 vccd1 vccd1 _8613__29/HI _8708_/A sky130_fd_sc_hd__conb_1
XFILLER_28_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7912_ _8099_/A _7978_/B vssd1 vssd1 vccd1 vccd1 _7913_/A sky130_fd_sc_hd__or2_1
XFILLER_36_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7843_ _7951_/A _7950_/A vssd1 vssd1 vccd1 vccd1 _7886_/A sky130_fd_sc_hd__nor2_2
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4986_ _5090_/A _5095_/C vssd1 vssd1 vccd1 vccd1 _5092_/A sky130_fd_sc_hd__or2_1
X_7774_ _7802_/A _7802_/B vssd1 vssd1 vccd1 vccd1 _7818_/B sky130_fd_sc_hd__xnor2_1
X_6725_ _6725_/A _6725_/B _6725_/C vssd1 vssd1 vccd1 vccd1 _6937_/A sky130_fd_sc_hd__or3_1
X_6656_ _7007_/A _6654_/Y _6680_/A vssd1 vssd1 vccd1 vccd1 _6657_/B sky130_fd_sc_hd__a21oi_2
X_6587_ _6829_/A vssd1 vssd1 vccd1 vccd1 _6812_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5607_ _5607_/A _5764_/B _5764_/C vssd1 vssd1 vccd1 vccd1 _5628_/A sky130_fd_sc_hd__or3_1
XFILLER_11_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8326_ _8326_/A _8326_/B _8326_/C vssd1 vssd1 vccd1 vccd1 _8326_/X sky130_fd_sc_hd__or3_1
X_5538_ _5538_/A _5538_/B _5427_/Y vssd1 vssd1 vccd1 vccd1 _5539_/B sky130_fd_sc_hd__or3b_1
X_8257_ _8257_/A _8257_/B vssd1 vssd1 vccd1 vccd1 _8285_/A sky130_fd_sc_hd__xnor2_1
XFILLER_3_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7208_ _7208_/A _7208_/B vssd1 vssd1 vccd1 vccd1 _7219_/B sky130_fd_sc_hd__xnor2_1
X_5469_ _5492_/B _5724_/A vssd1 vssd1 vccd1 vccd1 _6137_/A sky130_fd_sc_hd__xnor2_2
X_8188_ _8188_/A _8188_/B vssd1 vssd1 vccd1 vccd1 _8201_/C sky130_fd_sc_hd__xor2_1
X_7139_ _7139_/A _7132_/B vssd1 vssd1 vccd1 vccd1 _7139_/X sky130_fd_sc_hd__or2b_1
XFILLER_36_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8679__95 vssd1 vssd1 vccd1 vccd1 _8679__95/HI _8788_/A sky130_fd_sc_hd__conb_1
XFILLER_10_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4840_ _4840_/A vssd1 vssd1 vccd1 vccd1 _5031_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4771_ _4790_/A _4779_/A _4790_/B vssd1 vssd1 vccd1 vccd1 _4771_/X sky130_fd_sc_hd__or3_1
X_6510_ _7410_/A _7613_/B vssd1 vssd1 vccd1 vccd1 _6512_/A sky130_fd_sc_hd__and2_1
XFILLER_20_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7490_ _7766_/A _7489_/Y _4510_/A vssd1 vssd1 vccd1 vccd1 _7490_/Y sky130_fd_sc_hd__o21ai_1
X_6441_ _6433_/A _6445_/B _6434_/Y vssd1 vssd1 vccd1 vccd1 _6442_/B sky130_fd_sc_hd__a21o_1
XFILLER_9_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6372_ _6371_/B _8539_/Q _6366_/B _8541_/Q vssd1 vssd1 vccd1 vccd1 _6373_/C sky130_fd_sc_hd__a31o_1
X_5323_ _5359_/B _5322_/X vssd1 vssd1 vccd1 vccd1 _5323_/X sky130_fd_sc_hd__or2b_1
X_8111_ _8111_/A _8111_/B _8111_/C vssd1 vssd1 vccd1 vccd1 _8112_/B sky130_fd_sc_hd__nand3_1
X_5254_ _8493_/Q _5252_/A _5241_/X vssd1 vssd1 vccd1 vccd1 _5255_/B sky130_fd_sc_hd__o21ai_1
X_8042_ _8306_/A _8025_/X _7980_/Y vssd1 vssd1 vccd1 vccd1 _8044_/B sky130_fd_sc_hd__a21o_1
X_5185_ _5185_/A _5185_/B vssd1 vssd1 vccd1 vccd1 _5185_/Y sky130_fd_sc_hd__nand2_1
XFILLER_95_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7826_ _7697_/A _8305_/S _8113_/A vssd1 vssd1 vccd1 vccd1 _7826_/Y sky130_fd_sc_hd__o21ai_1
X_4969_ _4969_/A _4969_/B vssd1 vssd1 vccd1 vccd1 _5035_/D sky130_fd_sc_hd__or2_2
XFILLER_11_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7757_ _7756_/A _7756_/B _7837_/A _7755_/X vssd1 vssd1 vccd1 vccd1 _7758_/C sky130_fd_sc_hd__a2bb2o_1
X_6708_ _7079_/A _6708_/B vssd1 vssd1 vccd1 vccd1 _6731_/B sky130_fd_sc_hd__xnor2_1
XFILLER_22_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7688_ _7756_/A _7954_/A _7702_/A _7702_/B vssd1 vssd1 vccd1 vccd1 _7690_/B sky130_fd_sc_hd__o22a_1
X_6639_ _7033_/A vssd1 vssd1 vccd1 vccd1 _7175_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_22_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8309_ _8309_/A _8309_/B vssd1 vssd1 vccd1 vccd1 _8310_/B sky130_fd_sc_hd__xnor2_1
XFILLER_78_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6990_ _6990_/A _6990_/B vssd1 vssd1 vccd1 vccd1 _6991_/B sky130_fd_sc_hd__or2_1
XFILLER_92_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5941_ _5624_/C _5942_/B _5827_/B _5940_/Y vssd1 vssd1 vccd1 vccd1 _6015_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_61_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5872_ _5872_/A _5872_/B vssd1 vssd1 vccd1 vccd1 _5896_/B sky130_fd_sc_hd__xor2_1
X_4823_ _5087_/A _5112_/B vssd1 vssd1 vccd1 vccd1 _5090_/B sky130_fd_sc_hd__or2_1
X_7611_ _7731_/A _7885_/A vssd1 vssd1 vccd1 vccd1 _7621_/A sky130_fd_sc_hd__nor2_1
X_4754_ _4675_/B _4754_/B _4759_/A vssd1 vssd1 vccd1 vccd1 _4908_/A sky130_fd_sc_hd__and3b_1
XFILLER_21_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7542_ _7542_/A _7542_/B vssd1 vssd1 vccd1 vccd1 _7649_/B sky130_fd_sc_hd__and2_2
X_7473_ _8573_/Q vssd1 vssd1 vccd1 vccd1 _7507_/A sky130_fd_sc_hd__inv_2
X_4685_ _5370_/A _4685_/B _4690_/B vssd1 vssd1 vccd1 vccd1 _4686_/A sky130_fd_sc_hd__and3_1
X_6424_ _6455_/A _6424_/B _6424_/C vssd1 vssd1 vccd1 vccd1 _6424_/X sky130_fd_sc_hd__or3_1
X_6355_ _8535_/Q _6357_/C _6348_/X vssd1 vssd1 vccd1 vccd1 _6356_/B sky130_fd_sc_hd__o21ai_1
XFILLER_88_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6286_ _6293_/B _6286_/B vssd1 vssd1 vccd1 vccd1 _6289_/C sky130_fd_sc_hd__and2b_1
X_5306_ _8526_/Q _5322_/C _5300_/X _5305_/X vssd1 vssd1 vccd1 vccd1 _5306_/X sky130_fd_sc_hd__o31a_1
XFILLER_88_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5237_ _8487_/Q _8486_/Q _8488_/Q vssd1 vssd1 vccd1 vccd1 _5238_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8025_ _8025_/A _8249_/B vssd1 vssd1 vccd1 vccd1 _8025_/X sky130_fd_sc_hd__or2_1
XFILLER_84_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5168_ _4873_/A _5093_/B _5167_/X vssd1 vssd1 vccd1 vccd1 _5169_/C sky130_fd_sc_hd__o21ba_1
X_5099_ _5099_/A _5099_/B _5099_/C vssd1 vssd1 vccd1 vccd1 _5099_/X sky130_fd_sc_hd__or3_1
XFILLER_83_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8789_ _8789_/A _4385_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[36] sky130_fd_sc_hd__ebufn_8
XFILLER_52_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7809_ _8176_/A _7810_/B _7830_/B vssd1 vssd1 vccd1 vccd1 _7930_/A sky130_fd_sc_hd__o21ai_1
XFILLER_4_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8649__65 vssd1 vssd1 vccd1 vccd1 _8649__65/HI _8758_/A sky130_fd_sc_hd__conb_1
XFILLER_79_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4470_ _4470_/A _4470_/B _4470_/C _4470_/D vssd1 vssd1 vccd1 vccd1 _4495_/B sky130_fd_sc_hd__and4_2
XFILLER_7_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6140_ _6140_/A _6198_/B vssd1 vssd1 vccd1 vccd1 _6141_/B sky130_fd_sc_hd__xnor2_1
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6071_ _6071_/A _6071_/B vssd1 vssd1 vccd1 vccd1 _6073_/B sky130_fd_sc_hd__xnor2_1
X_5022_ _5035_/D _5022_/B _5022_/C _5022_/D vssd1 vssd1 vccd1 vccd1 _5022_/X sky130_fd_sc_hd__or4_1
XFILLER_78_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6973_ _7038_/A _7032_/C vssd1 vssd1 vccd1 vccd1 _7176_/B sky130_fd_sc_hd__nor2_1
X_8712_ _8712_/A _4294_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[29] sky130_fd_sc_hd__ebufn_8
X_5924_ _5924_/A _5924_/B vssd1 vssd1 vccd1 vccd1 _5957_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5855_ _5855_/A _5855_/B vssd1 vssd1 vccd1 vccd1 _5901_/A sky130_fd_sc_hd__or2_1
XFILLER_34_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4806_ _4921_/B _4886_/C vssd1 vssd1 vccd1 vccd1 _4993_/A sky130_fd_sc_hd__or2_2
XFILLER_21_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8574_ input3/X _8574_/D vssd1 vssd1 vccd1 vccd1 _8574_/Q sky130_fd_sc_hd__dfxtp_1
X_5786_ _5785_/Y _5754_/X _5932_/B vssd1 vssd1 vccd1 vccd1 _5868_/A sky130_fd_sc_hd__a21oi_4
X_4737_ _4737_/A _4738_/B vssd1 vssd1 vccd1 vccd1 _4755_/A sky130_fd_sc_hd__nor2_1
X_7525_ _7528_/B vssd1 vssd1 vccd1 vccd1 _7695_/B sky130_fd_sc_hd__clkbuf_2
X_4668_ _8419_/A vssd1 vssd1 vccd1 vccd1 _4668_/X sky130_fd_sc_hd__clkbuf_2
X_7456_ _8403_/A _7456_/B vssd1 vssd1 vccd1 vccd1 _7457_/A sky130_fd_sc_hd__and2_1
X_6407_ _7384_/B _7380_/A _8561_/Q _7391_/A vssd1 vssd1 vccd1 vccd1 _6407_/X sky130_fd_sc_hd__a31o_1
X_4599_ _4659_/A _4659_/B _5179_/B _4659_/D vssd1 vssd1 vccd1 vccd1 _4671_/B sky130_fd_sc_hd__nor4_2
X_7387_ _7377_/S _7382_/B _7381_/A vssd1 vssd1 vccd1 vccd1 _7388_/B sky130_fd_sc_hd__o21ai_1
X_6338_ _8530_/Q _6338_/B vssd1 vssd1 vccd1 vccd1 _6339_/B sky130_fd_sc_hd__or2_1
XFILLER_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6269_ _8507_/Q _6270_/A vssd1 vssd1 vccd1 vccd1 _6271_/A sky130_fd_sc_hd__or2b_1
XFILLER_88_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8008_ _8037_/B _8008_/B vssd1 vssd1 vccd1 vccd1 _8010_/B sky130_fd_sc_hd__xnor2_1
XFILLER_29_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5640_ _5718_/B _5639_/C _5639_/A vssd1 vssd1 vccd1 vccd1 _5669_/B sky130_fd_sc_hd__a21o_1
X_5571_ _5839_/A _6188_/B _5570_/X _5466_/A _5466_/Y vssd1 vssd1 vccd1 vccd1 _5586_/B
+ sky130_fd_sc_hd__a221o_1
X_7310_ _6792_/B _6792_/C _7310_/S vssd1 vssd1 vccd1 vccd1 _7312_/A sky130_fd_sc_hd__mux2_1
X_8290_ _8295_/A _8290_/B vssd1 vssd1 vccd1 vccd1 _8291_/B sky130_fd_sc_hd__xnor2_2
X_4522_ _8436_/Q _4527_/C vssd1 vssd1 vccd1 vccd1 _4526_/A sky130_fd_sc_hd__and2_1
X_4453_ _5104_/A vssd1 vssd1 vccd1 vccd1 _5099_/A sky130_fd_sc_hd__clkbuf_2
X_7241_ _7241_/A _7241_/B _7241_/C vssd1 vssd1 vccd1 vccd1 _7243_/A sky130_fd_sc_hd__and3_1
X_7172_ _7172_/A _7172_/B vssd1 vssd1 vccd1 vccd1 _7200_/A sky130_fd_sc_hd__xnor2_1
X_4384_ _4387_/A vssd1 vssd1 vccd1 vccd1 _4384_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6123_ _6044_/A _6043_/B _6043_/A vssd1 vssd1 vccd1 vccd1 _6223_/A sky130_fd_sc_hd__o21ba_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6054_ _5715_/A _6053_/Y _5685_/C _5661_/B vssd1 vssd1 vccd1 vccd1 _6075_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5005_ _5136_/C _5002_/X _5004_/X _4862_/A vssd1 vssd1 vccd1 vccd1 _5006_/D sky130_fd_sc_hd__o211a_1
XFILLER_85_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6956_ _6954_/A _6954_/Y _6910_/B _6955_/Y vssd1 vssd1 vccd1 vccd1 _6961_/A sky130_fd_sc_hd__o211ai_1
X_5907_ _5970_/A _5970_/B vssd1 vssd1 vccd1 vccd1 _5908_/B sky130_fd_sc_hd__xor2_1
X_6887_ _6871_/B _6884_/X _6878_/X _6883_/X vssd1 vssd1 vccd1 vccd1 _6888_/C sky130_fd_sc_hd__a211oi_1
XFILLER_22_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5838_ _5838_/A vssd1 vssd1 vccd1 vccd1 _6137_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_8557_ input3/X _8557_/D vssd1 vssd1 vccd1 vccd1 _8557_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5769_ _5776_/A _5776_/B _5823_/B vssd1 vssd1 vccd1 vccd1 _5824_/B sky130_fd_sc_hd__and3_1
X_7508_ _7508_/A _7507_/X vssd1 vssd1 vccd1 vccd1 _7680_/B sky130_fd_sc_hd__nor2b_2
X_8488_ input3/X _8488_/D vssd1 vssd1 vccd1 vccd1 _8488_/Q sky130_fd_sc_hd__dfxtp_1
X_7439_ _8574_/Q vssd1 vssd1 vccd1 vccd1 _7518_/A sky130_fd_sc_hd__inv_2
X_8619__35 vssd1 vssd1 vccd1 vccd1 _8619__35/HI _8714_/A sky130_fd_sc_hd__conb_1
XFILLER_49_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6810_ _6810_/A _6810_/B _6832_/C vssd1 vssd1 vccd1 vccd1 _7296_/B sky130_fd_sc_hd__and3_1
XFILLER_51_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7790_ _7638_/A _7672_/B _7788_/X _7789_/Y vssd1 vssd1 vccd1 vccd1 _7792_/B sky130_fd_sc_hd__a211oi_2
X_6741_ _6802_/B _6802_/C _6740_/A vssd1 vssd1 vccd1 vccd1 _6742_/C sky130_fd_sc_hd__a21o_1
XFILLER_50_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6672_ _6672_/A vssd1 vssd1 vccd1 vccd1 _7068_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_31_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5623_ _5721_/B _5622_/C _5622_/A vssd1 vssd1 vccd1 vccd1 _5633_/B sky130_fd_sc_hd__a21oi_1
X_8411_ _8412_/B _8428_/A vssd1 vssd1 vccd1 vccd1 _8421_/A sky130_fd_sc_hd__and2b_1
X_8342_ _8342_/A _8342_/B vssd1 vssd1 vccd1 vccd1 _8343_/B sky130_fd_sc_hd__xnor2_1
X_5554_ _5554_/A _5554_/B vssd1 vssd1 vccd1 vccd1 _5555_/C sky130_fd_sc_hd__or2_1
X_8273_ _8273_/A vssd1 vssd1 vccd1 vccd1 _8273_/Y sky130_fd_sc_hd__inv_2
X_5485_ _5485_/A _5485_/B vssd1 vssd1 vccd1 vccd1 _5609_/C sky130_fd_sc_hd__xor2_2
X_4505_ _8449_/Q _8452_/Q _8451_/Q vssd1 vssd1 vccd1 vccd1 _4506_/D sky130_fd_sc_hd__or3_1
X_7224_ _7234_/A _7234_/B vssd1 vssd1 vccd1 vccd1 _7226_/B sky130_fd_sc_hd__or2b_1
X_4436_ _4670_/A _4670_/B vssd1 vssd1 vccd1 vccd1 _4671_/A sky130_fd_sc_hd__or2_1
X_7155_ _7155_/A _7155_/B _7155_/C vssd1 vssd1 vccd1 vccd1 _7177_/A sky130_fd_sc_hd__nand3_2
X_4367_ _4369_/A vssd1 vssd1 vccd1 vccd1 _4367_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6106_ _6106_/A _6106_/B vssd1 vssd1 vccd1 vccd1 _6112_/A sky130_fd_sc_hd__nand2_1
X_4298_ _4301_/A vssd1 vssd1 vccd1 vccd1 _4298_/Y sky130_fd_sc_hd__inv_2
X_7086_ _7081_/A _7081_/B _7085_/Y vssd1 vssd1 vccd1 vccd1 _7143_/B sky130_fd_sc_hd__o21a_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6037_ _5952_/A _6037_/B vssd1 vssd1 vccd1 vccd1 _6037_/X sky130_fd_sc_hd__and2b_1
XFILLER_27_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7988_ _7989_/A _8252_/A vssd1 vssd1 vccd1 vccd1 _8047_/A sky130_fd_sc_hd__nand2_2
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6939_ _6939_/A _6939_/B _7323_/B vssd1 vssd1 vccd1 vccd1 _6940_/A sky130_fd_sc_hd__or3_1
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5270_ _8498_/Q _6392_/C _5270_/C vssd1 vssd1 vccd1 vccd1 _5277_/C sky130_fd_sc_hd__and3_1
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7911_ _7697_/A _8305_/S _7827_/X vssd1 vssd1 vccd1 vccd1 _7915_/A sky130_fd_sc_hd__o21a_1
XFILLER_36_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7842_ _7888_/B vssd1 vssd1 vccd1 vccd1 _7950_/A sky130_fd_sc_hd__buf_2
X_4985_ _4985_/A _5147_/B vssd1 vssd1 vccd1 vccd1 _5095_/C sky130_fd_sc_hd__or2_1
X_7773_ _7778_/A _7804_/C vssd1 vssd1 vccd1 vccd1 _7802_/B sky130_fd_sc_hd__xnor2_1
X_6724_ _6725_/A _6725_/C _6725_/B vssd1 vssd1 vccd1 vccd1 _6937_/C sky130_fd_sc_hd__o21ai_1
XFILLER_51_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6655_ _6655_/A vssd1 vssd1 vccd1 vccd1 _6680_/A sky130_fd_sc_hd__clkbuf_2
X_6586_ _6586_/A vssd1 vssd1 vccd1 vccd1 _6829_/A sky130_fd_sc_hd__clkbuf_2
X_5606_ _5488_/Y _5502_/A _5490_/B _5625_/A vssd1 vssd1 vccd1 vccd1 _5612_/A sky130_fd_sc_hd__a22o_1
X_8325_ _8326_/C _8275_/B _7854_/B _8274_/S vssd1 vssd1 vccd1 vccd1 _8325_/X sky130_fd_sc_hd__a2bb2o_1
X_5537_ _5685_/A _5537_/B vssd1 vssd1 vccd1 vccd1 _5538_/B sky130_fd_sc_hd__nor2_1
X_8256_ _8254_/X _8256_/B vssd1 vssd1 vccd1 vccd1 _8257_/B sky130_fd_sc_hd__and2b_1
XFILLER_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7207_ _7176_/B _7206_/B _7206_/X vssd1 vssd1 vccd1 vccd1 _7208_/B sky130_fd_sc_hd__a21bo_1
X_5468_ _5488_/A vssd1 vssd1 vccd1 vccd1 _5724_/A sky130_fd_sc_hd__clkbuf_2
X_4419_ _5380_/B vssd1 vssd1 vccd1 vccd1 _4715_/A sky130_fd_sc_hd__clkbuf_1
X_5399_ _5397_/X _5422_/A vssd1 vssd1 vccd1 vccd1 _5400_/B sky130_fd_sc_hd__and2b_1
X_8187_ _8198_/A _8198_/B _8199_/B vssd1 vssd1 vccd1 vccd1 _8201_/B sky130_fd_sc_hd__and3_1
X_7138_ _7138_/A _7138_/B vssd1 vssd1 vccd1 vccd1 _7165_/B sky130_fd_sc_hd__xnor2_1
XFILLER_59_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7069_ _7069_/A _7069_/B vssd1 vssd1 vccd1 vccd1 _7070_/B sky130_fd_sc_hd__nor2_1
XFILLER_14_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4770_ _4908_/B _4812_/A _4760_/Y _4929_/A vssd1 vssd1 vccd1 vccd1 _4909_/B sky130_fd_sc_hd__a211o_1
XFILLER_60_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6440_ _6440_/A _6440_/B vssd1 vssd1 vccd1 vccd1 _6442_/A sky130_fd_sc_hd__nor2_1
X_6371_ _8541_/Q _6371_/B _6371_/C vssd1 vssd1 vccd1 vccd1 _6375_/B sky130_fd_sc_hd__and3_1
X_8110_ _8111_/A _8111_/B _8111_/C vssd1 vssd1 vccd1 vccd1 _8110_/Y sky130_fd_sc_hd__a21oi_1
X_5322_ _5360_/A _5366_/A _5322_/C _5322_/D vssd1 vssd1 vccd1 vccd1 _5322_/X sky130_fd_sc_hd__or4_1
X_5253_ _8493_/Q _8492_/Q _5253_/C vssd1 vssd1 vccd1 vccd1 _5258_/C sky130_fd_sc_hd__and3_1
X_8041_ _8041_/A _8113_/A _8041_/C vssd1 vssd1 vccd1 vccd1 _8127_/A sky130_fd_sc_hd__and3_1
X_5184_ _4438_/A _4464_/B _4495_/B _5182_/Y _5183_/X vssd1 vssd1 vccd1 vccd1 _5185_/B
+ sky130_fd_sc_hd__o2111a_1
XFILLER_3_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7825_ _7825_/A vssd1 vssd1 vccd1 vccd1 _8113_/A sky130_fd_sc_hd__buf_2
X_4968_ _4968_/A _5117_/B _4945_/B vssd1 vssd1 vccd1 vccd1 _4972_/A sky130_fd_sc_hd__or3b_1
X_7756_ _7756_/A _7756_/B _7837_/A _7755_/X vssd1 vssd1 vccd1 vccd1 _7837_/B sky130_fd_sc_hd__or4bb_1
X_4899_ _4899_/A _4899_/B vssd1 vssd1 vccd1 vccd1 _5041_/C sky130_fd_sc_hd__nor2_2
X_6707_ _6796_/A _6796_/B vssd1 vssd1 vccd1 vccd1 _6708_/B sky130_fd_sc_hd__xor2_1
X_7687_ _7961_/A _8317_/B _7686_/X _7756_/A _7581_/Y vssd1 vssd1 vccd1 vccd1 _7702_/B
+ sky130_fd_sc_hd__a221o_1
X_6638_ _6733_/B _6645_/C _6645_/A vssd1 vssd1 vccd1 vccd1 _6896_/B sky130_fd_sc_hd__a21o_1
XFILLER_22_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6569_ _6569_/A _6569_/B vssd1 vssd1 vccd1 vccd1 _6819_/A sky130_fd_sc_hd__or2_2
X_8308_ _8308_/A _8308_/B vssd1 vssd1 vccd1 vccd1 _8309_/B sky130_fd_sc_hd__xnor2_1
XFILLER_3_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8239_ _8108_/A _8108_/B _8238_/X vssd1 vssd1 vccd1 vccd1 _8240_/B sky130_fd_sc_hd__a21oi_1
XFILLER_86_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5940_ _5940_/A vssd1 vssd1 vccd1 vccd1 _5940_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_18_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5871_ _5871_/A _5871_/B vssd1 vssd1 vccd1 vccd1 _5872_/B sky130_fd_sc_hd__and2_1
XFILLER_21_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7610_ _7635_/C _7720_/B vssd1 vssd1 vccd1 vccd1 _7623_/A sky130_fd_sc_hd__xnor2_1
XFILLER_33_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4822_ _4910_/A _4822_/B vssd1 vssd1 vccd1 vccd1 _5112_/B sky130_fd_sc_hd__or2_2
XFILLER_33_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4753_ _4822_/B vssd1 vssd1 vccd1 vccd1 _5138_/B sky130_fd_sc_hd__clkbuf_2
X_7541_ _7505_/A _7505_/B _7507_/X _7517_/X _7508_/A vssd1 vssd1 vccd1 vccd1 _7542_/B
+ sky130_fd_sc_hd__a311o_1
X_7472_ _7518_/A _7482_/B vssd1 vssd1 vccd1 vccd1 _7477_/B sky130_fd_sc_hd__or2_1
X_4684_ _4684_/A _4808_/A _4438_/A vssd1 vssd1 vccd1 vccd1 _4690_/B sky130_fd_sc_hd__or3b_1
X_6423_ _6439_/A _6433_/A _6445_/A vssd1 vssd1 vccd1 vccd1 _6424_/C sky130_fd_sc_hd__o21a_1
X_6354_ _8535_/Q _6357_/C vssd1 vssd1 vccd1 vccd1 _6356_/A sky130_fd_sc_hd__and2_1
X_6285_ _8523_/Q _5326_/B _6284_/X _5213_/X vssd1 vssd1 vccd1 vccd1 _8523_/D sky130_fd_sc_hd__o211a_1
X_5305_ _6274_/B _6270_/A _8520_/Q _5304_/Y vssd1 vssd1 vccd1 vccd1 _5305_/X sky130_fd_sc_hd__a31o_1
X_5236_ _8488_/Q _8487_/Q _8486_/Q vssd1 vssd1 vccd1 vccd1 _5240_/B sky130_fd_sc_hd__and3_1
X_8024_ _8024_/A vssd1 vssd1 vccd1 vccd1 _8249_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_84_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5167_ _4759_/A _4675_/B _4944_/B _5101_/S vssd1 vssd1 vccd1 vccd1 _5167_/X sky130_fd_sc_hd__o31a_1
XFILLER_68_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5098_ _4614_/A _5084_/X _5089_/X _5097_/X _5176_/S vssd1 vssd1 vccd1 vccd1 _5098_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_68_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8594__10 vssd1 vssd1 vccd1 vccd1 _8594__10/HI _8689_/A sky130_fd_sc_hd__conb_1
XFILLER_52_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8788_ _8788_/A _4384_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[35] sky130_fd_sc_hd__ebufn_8
XFILLER_12_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7808_ _7808_/A _8241_/A vssd1 vssd1 vccd1 vccd1 _7830_/B sky130_fd_sc_hd__xnor2_2
XFILLER_12_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7739_ _7840_/B _7738_/C _7738_/A vssd1 vssd1 vccd1 vccd1 _7752_/B sky130_fd_sc_hd__a21oi_1
XFILLER_33_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6070_ _5673_/B _6070_/B vssd1 vssd1 vccd1 vccd1 _6073_/A sky130_fd_sc_hd__and2b_1
XFILLER_85_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5021_ _5064_/C _5018_/X _5020_/X vssd1 vssd1 vccd1 vccd1 _5022_/D sky130_fd_sc_hd__o21a_1
XFILLER_66_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8711_ _8711_/A _4293_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[28] sky130_fd_sc_hd__ebufn_8
XFILLER_80_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6972_ _6972_/A vssd1 vssd1 vccd1 vccd1 _7038_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_53_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5923_ _5923_/A _5923_/B vssd1 vssd1 vccd1 vccd1 _5924_/B sky130_fd_sc_hd__xnor2_2
XFILLER_80_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5854_ _5916_/A _5854_/B vssd1 vssd1 vccd1 vccd1 _5872_/A sky130_fd_sc_hd__xnor2_1
X_4805_ _4805_/A _4809_/B vssd1 vssd1 vccd1 vccd1 _4886_/C sky130_fd_sc_hd__nor2_1
X_8573_ input3/X _8573_/D vssd1 vssd1 vccd1 vccd1 _8573_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5785_ _5785_/A _5785_/B vssd1 vssd1 vccd1 vccd1 _5785_/Y sky130_fd_sc_hd__nand2_1
X_7524_ _7537_/A _7524_/B vssd1 vssd1 vccd1 vccd1 _7528_/B sky130_fd_sc_hd__xor2_2
X_4736_ _4779_/A _4804_/A vssd1 vssd1 vccd1 vccd1 _5099_/C sky130_fd_sc_hd__nor2_2
XFILLER_21_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4667_ _4689_/A vssd1 vssd1 vccd1 vccd1 _8419_/A sky130_fd_sc_hd__buf_2
X_7455_ _7454_/Y _7452_/A _8430_/A vssd1 vssd1 vccd1 vccd1 _7456_/B sky130_fd_sc_hd__mux2_1
X_6406_ _6562_/B _7390_/A vssd1 vssd1 vccd1 vccd1 _7391_/A sky130_fd_sc_hd__or2b_1
X_7386_ _7386_/A _7386_/B vssd1 vssd1 vccd1 vccd1 _7388_/A sky130_fd_sc_hd__nor2_1
X_4598_ _5069_/A _4614_/A vssd1 vssd1 vccd1 vccd1 _4659_/D sky130_fd_sc_hd__nand2_1
X_6337_ _8530_/Q _6338_/B vssd1 vssd1 vccd1 vccd1 _6343_/C sky130_fd_sc_hd__and2_1
XFILLER_1_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6268_ _6268_/A vssd1 vssd1 vccd1 vccd1 _8520_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5219_ _8487_/Q _8486_/Q vssd1 vssd1 vccd1 vccd1 _6399_/A sky130_fd_sc_hd__or2_1
XFILLER_57_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6199_ _5851_/A _6141_/B _6198_/X vssd1 vssd1 vccd1 vccd1 _6200_/B sky130_fd_sc_hd__a21o_1
XFILLER_28_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8007_ _8007_/A _8037_/A vssd1 vssd1 vccd1 vccd1 _8008_/B sky130_fd_sc_hd__nor2_1
XFILLER_28_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5570_ _5839_/A _5846_/A vssd1 vssd1 vccd1 vccd1 _5570_/X sky130_fd_sc_hd__or2b_1
X_4521_ _4521_/A vssd1 vssd1 vccd1 vccd1 _8435_/D sky130_fd_sc_hd__clkbuf_1
X_4452_ _8454_/Q vssd1 vssd1 vccd1 vccd1 _5104_/A sky130_fd_sc_hd__clkbuf_2
X_7240_ _7240_/A vssd1 vssd1 vccd1 vccd1 _7241_/C sky130_fd_sc_hd__inv_2
X_7171_ _7171_/A _7171_/B vssd1 vssd1 vccd1 vccd1 _7338_/A sky130_fd_sc_hd__and2_1
X_4383_ _4387_/A vssd1 vssd1 vccd1 vccd1 _4383_/Y sky130_fd_sc_hd__inv_2
X_6122_ _6122_/A _6122_/B vssd1 vssd1 vccd1 vccd1 _6224_/A sky130_fd_sc_hd__xnor2_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6053_ _6053_/A _6053_/B vssd1 vssd1 vccd1 vccd1 _6053_/Y sky130_fd_sc_hd__nor2_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5004_ _5136_/A _5090_/B _5004_/C _5004_/D vssd1 vssd1 vccd1 vccd1 _5004_/X sky130_fd_sc_hd__or4_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6955_ _6909_/A _6909_/C _6909_/B vssd1 vssd1 vccd1 vccd1 _6955_/Y sky130_fd_sc_hd__o21ai_1
X_5906_ _5861_/A _5860_/B _5859_/B _5863_/A _5863_/B vssd1 vssd1 vccd1 vccd1 _5970_/B
+ sky130_fd_sc_hd__a32o_1
X_6886_ _6886_/A _6886_/B vssd1 vssd1 vccd1 vccd1 _6888_/B sky130_fd_sc_hd__xnor2_1
XFILLER_22_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5837_ _6188_/A _5940_/A vssd1 vssd1 vccd1 vccd1 _5927_/A sky130_fd_sc_hd__or2_1
X_8556_ input3/X _8556_/D vssd1 vssd1 vccd1 vccd1 _8556_/Q sky130_fd_sc_hd__dfxtp_1
X_5768_ _5767_/X _5725_/X _5724_/Y _5619_/A vssd1 vssd1 vccd1 vccd1 _5823_/B sky130_fd_sc_hd__a2bb2o_1
X_4719_ _4809_/B _4875_/B vssd1 vssd1 vccd1 vccd1 _5011_/A sky130_fd_sc_hd__nor2_1
X_8487_ input3/X _8487_/D vssd1 vssd1 vccd1 vccd1 _8487_/Q sky130_fd_sc_hd__dfxtp_1
X_7507_ _7507_/A _8470_/Q vssd1 vssd1 vccd1 vccd1 _7507_/X sky130_fd_sc_hd__or2_1
X_5699_ _5699_/A _5699_/B vssd1 vssd1 vccd1 vccd1 _5699_/X sky130_fd_sc_hd__or2_1
XFILLER_30_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7438_ _7459_/A _7438_/B vssd1 vssd1 vccd1 vccd1 _7438_/Y sky130_fd_sc_hd__nand2_1
X_7369_ _7372_/B _7372_/C vssd1 vssd1 vccd1 vccd1 _7369_/X sky130_fd_sc_hd__and2_1
XFILLER_89_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6740_ _6740_/A _6802_/B _6802_/C vssd1 vssd1 vccd1 vccd1 _6816_/A sky130_fd_sc_hd__nand3_1
XFILLER_90_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6671_ _6680_/A _6784_/A vssd1 vssd1 vccd1 vccd1 _6780_/A sky130_fd_sc_hd__nor2_2
X_5622_ _5622_/A _5721_/B _5622_/C vssd1 vssd1 vccd1 vccd1 _5633_/A sky130_fd_sc_hd__and3_1
X_8410_ _8410_/A _8410_/B vssd1 vssd1 vccd1 vccd1 _8584_/D sky130_fd_sc_hd__nor2_1
X_8341_ _8341_/A _8341_/B vssd1 vssd1 vccd1 vccd1 _8342_/B sky130_fd_sc_hd__xnor2_1
X_5553_ _5554_/A _5554_/B vssd1 vssd1 vccd1 vccd1 _5555_/B sky130_fd_sc_hd__nand2_1
X_4504_ _8448_/Q _8447_/Q _8450_/Q _8453_/Q vssd1 vssd1 vccd1 vccd1 _4506_/C sky130_fd_sc_hd__or4b_1
X_8272_ _8148_/A _8274_/S _8149_/B _8260_/C vssd1 vssd1 vccd1 vccd1 _8326_/C sky130_fd_sc_hd__a22oi_4
X_5484_ _5432_/B _5461_/A _5444_/B _5483_/Y vssd1 vssd1 vccd1 vccd1 _5485_/B sky130_fd_sc_hd__a31o_1
X_7223_ _7183_/A _7121_/A _7232_/A _7232_/B vssd1 vssd1 vccd1 vccd1 _7234_/B sky130_fd_sc_hd__a2bb2o_1
X_4435_ _4759_/A _4754_/B vssd1 vssd1 vccd1 vccd1 _4670_/B sky130_fd_sc_hd__nor2_1
XFILLER_6_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7154_ _7129_/A _7105_/C _7105_/A vssd1 vssd1 vccd1 vccd1 _7155_/C sky130_fd_sc_hd__a21o_1
X_4366_ _4369_/A vssd1 vssd1 vccd1 vccd1 _4366_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6105_ _6004_/A _6004_/B _6104_/Y vssd1 vssd1 vccd1 vccd1 _6211_/A sky130_fd_sc_hd__a21bo_1
X_4297_ _4301_/A vssd1 vssd1 vccd1 vccd1 _4297_/Y sky130_fd_sc_hd__inv_2
X_7085_ _7085_/A _7085_/B vssd1 vssd1 vccd1 vccd1 _7085_/Y sky130_fd_sc_hd__nand2_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6036_ _6036_/A _6036_/B vssd1 vssd1 vccd1 vccd1 _6160_/A sky130_fd_sc_hd__xnor2_1
XFILLER_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7987_ _8041_/A _8113_/A _8041_/C vssd1 vssd1 vccd1 vccd1 _8252_/A sky130_fd_sc_hd__nand3_2
X_6938_ _6938_/A _6938_/B vssd1 vssd1 vccd1 vccd1 _7009_/A sky130_fd_sc_hd__xnor2_1
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6869_ _7282_/A _6867_/C _6867_/B vssd1 vssd1 vccd1 vccd1 _6870_/D sky130_fd_sc_hd__a21o_1
XFILLER_22_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8539_ input3/X _8539_/D vssd1 vssd1 vccd1 vccd1 _8539_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7910_ _7939_/A _7939_/B vssd1 vssd1 vccd1 vccd1 _7935_/A sky130_fd_sc_hd__xnor2_1
XFILLER_48_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7841_ _7841_/A _7841_/B vssd1 vssd1 vccd1 vccd1 _7881_/A sky130_fd_sc_hd__nand2_1
XFILLER_63_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4984_ _5135_/B vssd1 vssd1 vccd1 vccd1 _5109_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_63_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7772_ _8176_/A _7772_/B vssd1 vssd1 vccd1 vccd1 _7804_/C sky130_fd_sc_hd__nor2_2
X_6723_ _6723_/A vssd1 vssd1 vccd1 vccd1 _6725_/B sky130_fd_sc_hd__inv_2
X_6654_ _6683_/A _6683_/B _7067_/B vssd1 vssd1 vccd1 vccd1 _6654_/Y sky130_fd_sc_hd__o21ai_1
X_5605_ _5504_/A _5504_/B _5604_/X vssd1 vssd1 vccd1 vccd1 _5622_/A sky130_fd_sc_hd__a21o_1
X_6585_ _6806_/A _6585_/B _6585_/C vssd1 vssd1 vccd1 vccd1 _6586_/A sky130_fd_sc_hd__and3b_1
XFILLER_11_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8324_ _8324_/A _8324_/B vssd1 vssd1 vccd1 vccd1 _8331_/A sky130_fd_sc_hd__xnor2_1
X_5536_ _5540_/A _5664_/B vssd1 vssd1 vccd1 vccd1 _5539_/A sky130_fd_sc_hd__xor2_1
X_8255_ _8255_/A _8255_/B _8255_/C vssd1 vssd1 vccd1 vccd1 _8256_/B sky130_fd_sc_hd__or3_1
X_5467_ _5467_/A vssd1 vssd1 vccd1 vccd1 _5488_/A sky130_fd_sc_hd__clkbuf_2
X_7206_ _7233_/B _7206_/B vssd1 vssd1 vccd1 vccd1 _7206_/X sky130_fd_sc_hd__or2_1
X_4418_ _8469_/Q vssd1 vssd1 vccd1 vccd1 _5380_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_59_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8186_ _8186_/A _8186_/B vssd1 vssd1 vccd1 vccd1 _8199_/B sky130_fd_sc_hd__xnor2_1
X_5398_ _7518_/B _8513_/Q vssd1 vssd1 vccd1 vccd1 _5422_/A sky130_fd_sc_hd__or2b_1
X_7137_ _7138_/A _7138_/B vssd1 vssd1 vccd1 vccd1 _7137_/X sky130_fd_sc_hd__and2_1
X_4349_ _4351_/A vssd1 vssd1 vccd1 vccd1 _4349_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7068_ _7202_/A _7068_/B vssd1 vssd1 vccd1 vccd1 _7070_/A sky130_fd_sc_hd__nor2_1
XFILLER_86_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6019_ _6019_/A _6019_/B vssd1 vssd1 vccd1 vccd1 _6020_/B sky130_fd_sc_hd__or2_1
XFILLER_54_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6370_ _6371_/B _6371_/C _6369_/Y vssd1 vssd1 vccd1 vccd1 _8540_/D sky130_fd_sc_hd__a21oi_1
X_5321_ _5339_/B _5335_/A _5345_/B vssd1 vssd1 vccd1 vccd1 _5322_/D sky130_fd_sc_hd__o21a_1
X_8040_ _7995_/A _7995_/B _8039_/X vssd1 vssd1 vccd1 vccd1 _8088_/A sky130_fd_sc_hd__a21boi_1
XFILLER_87_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5252_ _5252_/A _5252_/B vssd1 vssd1 vccd1 vccd1 _8492_/D sky130_fd_sc_hd__nor2_1
X_5183_ _5526_/B _4706_/A _4466_/B _4715_/A _4698_/A vssd1 vssd1 vccd1 vccd1 _5183_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7824_ _7824_/A _8105_/B vssd1 vssd1 vccd1 vccd1 _7825_/A sky130_fd_sc_hd__or2_1
X_4967_ _5010_/C vssd1 vssd1 vccd1 vccd1 _5117_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7755_ _7839_/B _7754_/C _7754_/A vssd1 vssd1 vccd1 vccd1 _7755_/X sky130_fd_sc_hd__a21o_1
X_4898_ _4898_/A _5171_/C _4938_/A vssd1 vssd1 vccd1 vccd1 _4906_/D sky130_fd_sc_hd__or3_1
X_6706_ _6727_/A _6727_/B _6705_/Y vssd1 vssd1 vccd1 vccd1 _6796_/B sky130_fd_sc_hd__a21oi_1
X_7686_ _7961_/A _7969_/A vssd1 vssd1 vccd1 vccd1 _7686_/X sky130_fd_sc_hd__or2b_1
X_6637_ _6892_/A _6990_/A vssd1 vssd1 vccd1 vccd1 _6645_/A sky130_fd_sc_hd__and2_1
X_6568_ _6714_/A _6784_/A _6655_/A vssd1 vssd1 vccd1 vccd1 _6569_/B sky130_fd_sc_hd__a21o_1
X_8307_ _8227_/Y _8306_/Y _8105_/B vssd1 vssd1 vccd1 vccd1 _8308_/B sky130_fd_sc_hd__a21o_1
X_5519_ _5520_/A _5520_/B vssd1 vssd1 vccd1 vccd1 _5521_/A sky130_fd_sc_hd__or2_1
X_6499_ _6499_/A _6499_/B vssd1 vssd1 vccd1 vccd1 _6500_/B sky130_fd_sc_hd__nor2_2
X_8238_ _8109_/B _8238_/B vssd1 vssd1 vccd1 vccd1 _8238_/X sky130_fd_sc_hd__and2b_1
XFILLER_78_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8169_ _8169_/A _8169_/B vssd1 vssd1 vccd1 vccd1 _8170_/B sky130_fd_sc_hd__xnor2_1
XFILLER_59_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5870_ _5870_/A _5870_/B vssd1 vssd1 vccd1 vccd1 _5871_/B sky130_fd_sc_hd__nand2_1
XFILLER_33_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4821_ _4938_/A _4871_/A vssd1 vssd1 vccd1 vccd1 _4910_/A sky130_fd_sc_hd__or2_1
X_4752_ _4855_/A _5074_/B vssd1 vssd1 vccd1 vccd1 _4822_/B sky130_fd_sc_hd__or2_1
X_7540_ _7540_/A _7539_/Y vssd1 vssd1 vccd1 vccd1 _7649_/A sky130_fd_sc_hd__nor2b_4
X_4683_ _5207_/A _4808_/A _4438_/A vssd1 vssd1 vccd1 vccd1 _4685_/B sky130_fd_sc_hd__o21bai_1
X_7471_ _8573_/Q _6348_/X _7470_/X vssd1 vssd1 vccd1 vccd1 _8573_/D sky130_fd_sc_hd__a21bo_1
X_6422_ _6541_/A _6419_/X _6452_/A _8556_/Q vssd1 vssd1 vccd1 vccd1 _6422_/Y sky130_fd_sc_hd__a31oi_1
X_6353_ _6357_/C _6353_/B vssd1 vssd1 vccd1 vccd1 _8534_/D sky130_fd_sc_hd__nor2_1
X_5304_ _6289_/A vssd1 vssd1 vccd1 vccd1 _5304_/Y sky130_fd_sc_hd__inv_2
X_6284_ _5304_/Y _6289_/B _6283_/Y _5368_/B vssd1 vssd1 vccd1 vccd1 _6284_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5235_ _5235_/A vssd1 vssd1 vccd1 vccd1 _8487_/D sky130_fd_sc_hd__clkbuf_1
X_8023_ _8023_/A _8023_/B vssd1 vssd1 vccd1 vccd1 _8341_/A sky130_fd_sc_hd__nand2_1
XFILLER_96_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5166_ _5151_/C _5159_/X _5160_/X _5165_/X _5156_/C vssd1 vssd1 vccd1 vccd1 _5166_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_68_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5097_ _5135_/B _5096_/X _4624_/A vssd1 vssd1 vccd1 vccd1 _5097_/X sky130_fd_sc_hd__o21a_1
XFILLER_56_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8787_ _8787_/A _4383_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[34] sky130_fd_sc_hd__ebufn_8
XFILLER_12_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5999_ _5999_/A _5999_/B vssd1 vssd1 vccd1 vccd1 _6000_/B sky130_fd_sc_hd__nor2_1
X_7807_ _7914_/A vssd1 vssd1 vccd1 vccd1 _8241_/A sky130_fd_sc_hd__buf_2
X_7738_ _7738_/A _7840_/B _7738_/C vssd1 vssd1 vccd1 vccd1 _7752_/A sky130_fd_sc_hd__and3_1
X_7669_ _7715_/A _7669_/B vssd1 vssd1 vccd1 vccd1 _7671_/B sky130_fd_sc_hd__and2_1
XFILLER_58_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5020_ _5136_/B _5020_/B _5020_/C _5020_/D vssd1 vssd1 vccd1 vccd1 _5020_/X sky130_fd_sc_hd__or4_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8710_ _8710_/A _4292_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[27] sky130_fd_sc_hd__ebufn_8
XFILLER_80_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6971_ _6971_/A _6971_/B vssd1 vssd1 vccd1 vccd1 _7035_/B sky130_fd_sc_hd__xnor2_2
XFILLER_19_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5922_ _6010_/A _5922_/B vssd1 vssd1 vccd1 vccd1 _5923_/B sky130_fd_sc_hd__nor2_2
X_5853_ _5853_/A _5853_/B vssd1 vssd1 vccd1 vccd1 _5854_/B sky130_fd_sc_hd__xor2_2
XFILLER_21_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4804_ _4804_/A _4818_/B vssd1 vssd1 vccd1 vccd1 _4921_/B sky130_fd_sc_hd__nor2_1
X_8572_ input3/X _8572_/D vssd1 vssd1 vccd1 vccd1 _8572_/Q sky130_fd_sc_hd__dfxtp_1
X_5784_ _6021_/A vssd1 vssd1 vccd1 vccd1 _5932_/B sky130_fd_sc_hd__buf_2
X_4735_ _4735_/A _4735_/B _4754_/B _4748_/D vssd1 vssd1 vccd1 vccd1 _4804_/A sky130_fd_sc_hd__or4b_2
X_7523_ _7921_/A vssd1 vssd1 vccd1 vccd1 _7813_/A sky130_fd_sc_hd__clkbuf_2
X_4666_ _4705_/A vssd1 vssd1 vccd1 vccd1 _4790_/A sky130_fd_sc_hd__buf_2
X_7454_ _8570_/Q _7454_/B vssd1 vssd1 vccd1 vccd1 _7454_/Y sky130_fd_sc_hd__xnor2_1
X_4597_ _4624_/A vssd1 vssd1 vccd1 vccd1 _5069_/A sky130_fd_sc_hd__clkbuf_2
X_6405_ _8564_/Q vssd1 vssd1 vccd1 vccd1 _6562_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_7385_ _7384_/B _7390_/A vssd1 vssd1 vccd1 vccd1 _7386_/B sky130_fd_sc_hd__and2b_1
X_6336_ _6336_/A vssd1 vssd1 vccd1 vccd1 _8529_/D sky130_fd_sc_hd__clkbuf_1
X_6267_ _5332_/A _5328_/A _6267_/S vssd1 vssd1 vccd1 vccd1 _6268_/A sky130_fd_sc_hd__mux2_1
X_5218_ _8560_/Q _5202_/A _5217_/X _5213_/X vssd1 vssd1 vccd1 vccd1 _8485_/D sky130_fd_sc_hd__o211a_1
X_8654__70 vssd1 vssd1 vccd1 vccd1 _8654__70/HI _8763_/A sky130_fd_sc_hd__conb_1
X_6198_ _6140_/A _6198_/B vssd1 vssd1 vccd1 vccd1 _6198_/X sky130_fd_sc_hd__and2b_1
X_8006_ _8367_/B _7808_/A _8113_/A vssd1 vssd1 vccd1 vccd1 _8007_/A sky130_fd_sc_hd__a21oi_1
X_5149_ _5173_/A _5149_/B vssd1 vssd1 vccd1 vccd1 _5156_/C sky130_fd_sc_hd__or2_1
XFILLER_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4520_ _4527_/C _4575_/A _4520_/C vssd1 vssd1 vccd1 vccd1 _4521_/A sky130_fd_sc_hd__and3b_1
X_4451_ _8455_/Q vssd1 vssd1 vccd1 vccd1 _5064_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7170_ _7345_/A _7345_/B _7345_/C vssd1 vssd1 vccd1 vccd1 _7171_/B sky130_fd_sc_hd__o21ai_1
X_4382_ _4382_/A vssd1 vssd1 vccd1 vccd1 _4387_/A sky130_fd_sc_hd__buf_2
X_6121_ _6121_/A vssd1 vssd1 vccd1 vccd1 _6122_/B sky130_fd_sc_hd__inv_2
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6052_ _6170_/A _6236_/B vssd1 vssd1 vccd1 vccd1 _6241_/A sky130_fd_sc_hd__xnor2_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5003_ _5092_/A _4987_/X _4873_/A vssd1 vssd1 vccd1 vccd1 _5004_/D sky130_fd_sc_hd__o21a_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6954_ _6954_/A _6954_/B _6954_/C vssd1 vssd1 vccd1 vccd1 _6954_/Y sky130_fd_sc_hd__nor3_2
XFILLER_53_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5905_ _6210_/A _5905_/B vssd1 vssd1 vccd1 vccd1 _5970_/A sky130_fd_sc_hd__xnor2_1
X_6885_ _6878_/X _6883_/X _6871_/B _6884_/X vssd1 vssd1 vccd1 vccd1 _6888_/A sky130_fd_sc_hd__o211a_1
XFILLER_14_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5836_ _5836_/A _5835_/X vssd1 vssd1 vccd1 vccd1 _5844_/A sky130_fd_sc_hd__or2b_1
XFILLER_22_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8555_ input3/X _8555_/D vssd1 vssd1 vccd1 vccd1 _8555_/Q sky130_fd_sc_hd__dfxtp_1
X_5767_ _5767_/A _5767_/B vssd1 vssd1 vccd1 vccd1 _5767_/X sky130_fd_sc_hd__or2_1
X_4718_ _4718_/A _4748_/B _4759_/B _4725_/A vssd1 vssd1 vccd1 vccd1 _4875_/B sky130_fd_sc_hd__or4b_4
X_8486_ input3/X _8486_/D vssd1 vssd1 vccd1 vccd1 _8486_/Q sky130_fd_sc_hd__dfxtp_1
X_5698_ _5698_/A _5698_/B vssd1 vssd1 vccd1 vccd1 _5747_/B sky130_fd_sc_hd__nand2_1
XFILLER_5_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7506_ _7507_/A _7506_/B vssd1 vssd1 vccd1 vccd1 _7508_/A sky130_fd_sc_hd__and2_1
X_4649_ _4711_/A _4649_/B vssd1 vssd1 vccd1 vccd1 _4656_/S sky130_fd_sc_hd__nand2_1
X_7437_ _7452_/A _8570_/Q _8573_/Q vssd1 vssd1 vccd1 vccd1 _7438_/B sky130_fd_sc_hd__a21oi_1
X_7368_ _7372_/B _7372_/C vssd1 vssd1 vccd1 vccd1 _7368_/Y sky130_fd_sc_hd__nor2_1
X_6319_ _8532_/Q _8538_/Q _8537_/Q _6319_/D vssd1 vssd1 vccd1 vccd1 _6320_/C sky130_fd_sc_hd__and4bb_1
X_7299_ _7299_/A _7299_/B vssd1 vssd1 vccd1 vccd1 _7300_/B sky130_fd_sc_hd__xnor2_1
XFILLER_39_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6670_ _6714_/B _6714_/C _6672_/A _7069_/B vssd1 vssd1 vccd1 vccd1 _6675_/A sky130_fd_sc_hd__or4_2
X_5621_ _5620_/A _5620_/B _5619_/X vssd1 vssd1 vccd1 vccd1 _5622_/C sky130_fd_sc_hd__o21bai_1
X_8340_ _8285_/A _8338_/X _8339_/X vssd1 vssd1 vccd1 vccd1 _8341_/B sky130_fd_sc_hd__o21a_1
X_5552_ _5599_/A _5552_/B vssd1 vssd1 vccd1 vccd1 _5554_/B sky130_fd_sc_hd__and2_1
X_8271_ _8159_/A _8159_/B _8270_/X vssd1 vssd1 vccd1 vccd1 _8334_/A sky130_fd_sc_hd__a21bo_1
X_4503_ _8436_/Q _8435_/Q _8438_/Q _8437_/Q vssd1 vssd1 vccd1 vccd1 _4506_/B sky130_fd_sc_hd__or4_1
X_5483_ _5497_/A vssd1 vssd1 vccd1 vccd1 _5483_/Y sky130_fd_sc_hd__inv_2
X_4434_ _4761_/B vssd1 vssd1 vccd1 vccd1 _4754_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_7222_ _7233_/A _6969_/A _7180_/B _7221_/X vssd1 vssd1 vccd1 vccd1 _7232_/B sky130_fd_sc_hd__o31a_1
XFILLER_6_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7153_ _7153_/A _7153_/B vssd1 vssd1 vccd1 vccd1 _7155_/B sky130_fd_sc_hd__and2_1
X_4365_ _4369_/A vssd1 vssd1 vccd1 vccd1 _4365_/Y sky130_fd_sc_hd__inv_2
X_7084_ _7065_/A _7082_/X _7083_/X _7019_/Y vssd1 vssd1 vccd1 vccd1 _7143_/A sky130_fd_sc_hd__o211a_1
XFILLER_58_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6104_ _6104_/A _6177_/A vssd1 vssd1 vccd1 vccd1 _6104_/Y sky130_fd_sc_hd__nand2_1
X_4296_ _4296_/A vssd1 vssd1 vccd1 vccd1 _4301_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_86_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8624__40 vssd1 vssd1 vccd1 vccd1 _8624__40/HI _8719_/A sky130_fd_sc_hd__conb_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6035_ _6154_/B _6147_/A vssd1 vssd1 vccd1 vccd1 _6036_/B sky130_fd_sc_hd__xnor2_1
XFILLER_86_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7986_ _7986_/A _7986_/B vssd1 vssd1 vccd1 vccd1 _7989_/A sky130_fd_sc_hd__xor2_1
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6937_ _6937_/A _6937_/B _6937_/C vssd1 vssd1 vccd1 vccd1 _6945_/A sky130_fd_sc_hd__nand3_1
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6868_ _6826_/A _6817_/B _6817_/C vssd1 vssd1 vccd1 vccd1 _6870_/C sky130_fd_sc_hd__a21o_1
X_5819_ _5814_/A _5814_/B _5818_/Y vssd1 vssd1 vccd1 vccd1 _5873_/A sky130_fd_sc_hd__o21a_1
X_8538_ input3/X _8538_/D vssd1 vssd1 vccd1 vccd1 _8538_/Q sky130_fd_sc_hd__dfxtp_1
X_6799_ _7176_/A _6810_/A vssd1 vssd1 vccd1 vccd1 _7291_/A sky130_fd_sc_hd__nor2_1
XFILLER_10_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8469_ input3/X _8469_/D vssd1 vssd1 vccd1 vccd1 _8469_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_49_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7840_ _7736_/A _7840_/B vssd1 vssd1 vccd1 vccd1 _7877_/B sky130_fd_sc_hd__and2b_1
XFILLER_91_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4983_ _5069_/A _5146_/A _4965_/X _4982_/X _4863_/X vssd1 vssd1 vccd1 vccd1 _4983_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_23_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7771_ _7528_/B _7921_/B _8023_/B vssd1 vssd1 vccd1 vccd1 _7772_/B sky130_fd_sc_hd__a21oi_1
X_6722_ _7054_/A _6926_/B vssd1 vssd1 vccd1 vccd1 _6723_/A sky130_fd_sc_hd__nor2_1
X_6653_ _6683_/A _7067_/B _6683_/B vssd1 vssd1 vccd1 vccd1 _7007_/A sky130_fd_sc_hd__or3_2
X_5604_ _5518_/C _5604_/B vssd1 vssd1 vccd1 vccd1 _5604_/X sky130_fd_sc_hd__and2b_1
X_6584_ _6584_/A _6632_/A vssd1 vssd1 vccd1 vccd1 _6585_/B sky130_fd_sc_hd__nand2_1
XFILLER_11_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8323_ _8323_/A _8323_/B vssd1 vssd1 vccd1 vccd1 _8324_/B sky130_fd_sc_hd__xnor2_1
X_5535_ _5541_/B _5535_/B vssd1 vssd1 vccd1 vccd1 _5664_/B sky130_fd_sc_hd__xnor2_2
X_8254_ _8255_/A _8255_/B _8255_/C vssd1 vssd1 vccd1 vccd1 _8254_/X sky130_fd_sc_hd__o21a_1
X_5466_ _5466_/A _5518_/C vssd1 vssd1 vccd1 vccd1 _5466_/Y sky130_fd_sc_hd__nor2_1
X_4417_ _4466_/B vssd1 vssd1 vccd1 vccd1 _4698_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_7205_ _7205_/A _7205_/B vssd1 vssd1 vccd1 vccd1 _7208_/A sky130_fd_sc_hd__nand2_1
X_5397_ _8513_/Q _8471_/Q vssd1 vssd1 vccd1 vccd1 _5397_/X sky130_fd_sc_hd__and2b_1
X_8185_ _8186_/A _8186_/B vssd1 vssd1 vccd1 vccd1 _8201_/A sky130_fd_sc_hd__and2b_1
X_7136_ _7136_/A _7136_/B vssd1 vssd1 vccd1 vccd1 _7138_/B sky130_fd_sc_hd__xor2_1
X_4348_ _4351_/A vssd1 vssd1 vccd1 vccd1 _4348_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4279_ _4283_/A vssd1 vssd1 vccd1 vccd1 _4279_/Y sky130_fd_sc_hd__inv_2
X_7067_ _7248_/A _7067_/B vssd1 vssd1 vccd1 vccd1 _7121_/A sky130_fd_sc_hd__nand2_2
XFILLER_74_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6018_ _6019_/A _6019_/B vssd1 vssd1 vccd1 vccd1 _6020_/A sky130_fd_sc_hd__nand2_1
XFILLER_39_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7969_ _7969_/A _8142_/A vssd1 vssd1 vccd1 vccd1 _8319_/A sky130_fd_sc_hd__nor2_1
XFILLER_42_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5320_ _5360_/B vssd1 vssd1 vccd1 vccd1 _5359_/B sky130_fd_sc_hd__clkbuf_1
X_5251_ _8492_/Q _5253_/C _5241_/X vssd1 vssd1 vccd1 vccd1 _5252_/B sky130_fd_sc_hd__o21ai_1
XFILLER_5_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5182_ _4639_/B _5178_/Y _4655_/X _5181_/X vssd1 vssd1 vccd1 vccd1 _5182_/Y sky130_fd_sc_hd__o31ai_1
XFILLER_95_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7823_ _7978_/B vssd1 vssd1 vccd1 vccd1 _8105_/B sky130_fd_sc_hd__clkbuf_2
X_7754_ _7754_/A _7839_/B _7754_/C vssd1 vssd1 vccd1 vccd1 _7837_/A sky130_fd_sc_hd__nand3_1
X_4966_ _4966_/A _4975_/C vssd1 vssd1 vccd1 vccd1 _5010_/C sky130_fd_sc_hd__or2_1
X_6705_ _6705_/A _6705_/B vssd1 vssd1 vccd1 vccd1 _6705_/Y sky130_fd_sc_hd__nor2_1
XFILLER_51_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4897_ _4897_/A vssd1 vssd1 vccd1 vccd1 _4898_/A sky130_fd_sc_hd__clkbuf_2
X_7685_ _7885_/A vssd1 vssd1 vccd1 vccd1 _7961_/A sky130_fd_sc_hd__buf_2
X_6636_ _6914_/C _6919_/A _6554_/Y vssd1 vssd1 vccd1 vccd1 _6990_/A sky130_fd_sc_hd__o21a_2
X_6567_ _6513_/X _6570_/B _6570_/C _6512_/A vssd1 vssd1 vccd1 vccd1 _6655_/A sky130_fd_sc_hd__a31o_1
XFILLER_3_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8306_ _8306_/A _8306_/B vssd1 vssd1 vccd1 vccd1 _8306_/Y sky130_fd_sc_hd__nand2_1
X_5518_ _6188_/A _5637_/A _5518_/C _5846_/A vssd1 vssd1 vccd1 vccd1 _5520_/B sky130_fd_sc_hd__or4b_2
X_6498_ _8469_/Q _8552_/Q vssd1 vssd1 vccd1 vccd1 _6499_/B sky130_fd_sc_hd__and2b_1
X_8237_ _8237_/A _8237_/B vssd1 vssd1 vccd1 vccd1 _8240_/A sky130_fd_sc_hd__xnor2_1
X_5449_ _5938_/A vssd1 vssd1 vccd1 vccd1 _6188_/A sky130_fd_sc_hd__clkbuf_2
X_8168_ _8168_/A _8221_/B vssd1 vssd1 vccd1 vccd1 _8169_/B sky130_fd_sc_hd__xnor2_1
X_7119_ _7202_/B _7148_/B _7116_/B vssd1 vssd1 vccd1 vccd1 _7126_/C sky130_fd_sc_hd__o21ai_1
XFILLER_74_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8099_ _8099_/A _8099_/B vssd1 vssd1 vccd1 vccd1 _8229_/A sky130_fd_sc_hd__or2_1
XFILLER_47_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4820_ _5080_/B _4906_/B vssd1 vssd1 vccd1 vccd1 _4871_/A sky130_fd_sc_hd__or2_1
XFILLER_61_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4751_ _4996_/A _4885_/A vssd1 vssd1 vccd1 vccd1 _5074_/B sky130_fd_sc_hd__or2_1
XFILLER_33_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4682_ _4689_/A vssd1 vssd1 vccd1 vccd1 _5370_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7470_ _7466_/X _7467_/X _7468_/Y _8426_/A vssd1 vssd1 vccd1 vccd1 _7470_/X sky130_fd_sc_hd__a211o_1
X_6421_ _6455_/A _6450_/B vssd1 vssd1 vccd1 vccd1 _6452_/A sky130_fd_sc_hd__or2_1
X_6352_ _8534_/Q _6350_/A _6331_/B vssd1 vssd1 vccd1 vccd1 _6353_/B sky130_fd_sc_hd__o21ai_1
X_6283_ _5304_/Y _6282_/B _6282_/A vssd1 vssd1 vccd1 vccd1 _6283_/Y sky130_fd_sc_hd__a21oi_1
X_5303_ _6281_/A _6281_/B vssd1 vssd1 vccd1 vccd1 _6289_/A sky130_fd_sc_hd__and2_1
XFILLER_69_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5234_ _6399_/A _5291_/A _5234_/C vssd1 vssd1 vccd1 vccd1 _5235_/A sky130_fd_sc_hd__and3_1
X_8022_ _8241_/A _8022_/B vssd1 vssd1 vccd1 vccd1 _8092_/A sky130_fd_sc_hd__nand2_1
X_5165_ _5059_/X _4921_/X _5159_/X _5164_/X vssd1 vssd1 vccd1 vccd1 _5165_/X sky130_fd_sc_hd__o31a_1
X_5096_ _4596_/A _5091_/X _5092_/X _5095_/X vssd1 vssd1 vccd1 vccd1 _5096_/X sky130_fd_sc_hd__o211a_1
XFILLER_83_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7806_ _7770_/A _8023_/B _7916_/A vssd1 vssd1 vccd1 vccd1 _7914_/A sky130_fd_sc_hd__mux2_2
X_8786_ _8786_/A _4381_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[33] sky130_fd_sc_hd__ebufn_8
X_5998_ _5999_/A _5999_/B vssd1 vssd1 vccd1 vccd1 _6110_/B sky130_fd_sc_hd__and2_1
XFILLER_33_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4949_ _4949_/A _4949_/B vssd1 vssd1 vccd1 vccd1 _4949_/Y sky130_fd_sc_hd__nand2_1
XFILLER_12_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7737_ _7736_/A _7736_/B _7735_/X vssd1 vssd1 vccd1 vccd1 _7738_/C sky130_fd_sc_hd__o21bai_1
XFILLER_20_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7668_ _7668_/A _7668_/B vssd1 vssd1 vccd1 vccd1 _7669_/B sky130_fd_sc_hd__nand2_1
X_6619_ _6618_/B _6618_/C _6804_/B vssd1 vssd1 vccd1 vccd1 _6620_/C sky130_fd_sc_hd__a21o_1
XFILLER_20_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7599_ _8462_/Q _8423_/A vssd1 vssd1 vccd1 vccd1 _7612_/A sky130_fd_sc_hd__or2b_1
XFILLER_94_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6970_ _7034_/S _6970_/B vssd1 vssd1 vccd1 vccd1 _6971_/B sky130_fd_sc_hd__xnor2_2
XFILLER_26_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5921_ _6006_/A _5921_/B vssd1 vssd1 vccd1 vccd1 _5922_/B sky130_fd_sc_hd__and2_1
XFILLER_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5852_ _5923_/A _5852_/B vssd1 vssd1 vccd1 vccd1 _5853_/B sky130_fd_sc_hd__nor2_1
X_4803_ _4747_/A _4750_/A _4786_/B vssd1 vssd1 vccd1 vccd1 _4993_/B sky130_fd_sc_hd__a21oi_1
XFILLER_61_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5783_ _5783_/A _5783_/B vssd1 vssd1 vccd1 vccd1 _5788_/A sky130_fd_sc_hd__xor2_2
X_8571_ input3/X _8571_/D vssd1 vssd1 vccd1 vccd1 _8571_/Q sky130_fd_sc_hd__dfxtp_1
X_4734_ _4767_/A vssd1 vssd1 vccd1 vccd1 _4779_/A sky130_fd_sc_hd__clkbuf_2
X_7522_ _7526_/B vssd1 vssd1 vccd1 vccd1 _7983_/A sky130_fd_sc_hd__clkbuf_2
X_4665_ _4748_/B _4766_/B vssd1 vssd1 vccd1 vccd1 _4705_/A sky130_fd_sc_hd__nand2_1
X_7453_ _7453_/A _7453_/B vssd1 vssd1 vccd1 vccd1 _7454_/B sky130_fd_sc_hd__nand2_1
X_4596_ _4596_/A vssd1 vssd1 vccd1 vccd1 _5179_/B sky130_fd_sc_hd__clkbuf_2
X_6404_ _8562_/Q vssd1 vssd1 vccd1 vccd1 _7380_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7384_ _7390_/A _7384_/B vssd1 vssd1 vccd1 vccd1 _7386_/A sky130_fd_sc_hd__and2b_1
X_6335_ _6338_/B _6335_/B _6389_/B vssd1 vssd1 vccd1 vccd1 _6336_/A sky130_fd_sc_hd__and3b_1
XFILLER_88_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8005_ _8003_/Y _8005_/B vssd1 vssd1 vccd1 vccd1 _8037_/B sky130_fd_sc_hd__and2b_1
X_6266_ _8520_/Q vssd1 vssd1 vccd1 vccd1 _6267_/S sky130_fd_sc_hd__inv_2
X_5217_ _8485_/Q _5217_/B vssd1 vssd1 vccd1 vccd1 _5217_/X sky130_fd_sc_hd__or2_1
XFILLER_69_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6197_ _6155_/A _6156_/A _6155_/B vssd1 vssd1 vccd1 vccd1 _6201_/A sky130_fd_sc_hd__o21ba_1
X_5148_ _5148_/A _5148_/B _5148_/C _5160_/D vssd1 vssd1 vccd1 vccd1 _5148_/X sky130_fd_sc_hd__or4_1
XFILLER_28_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5079_ _4938_/A _5074_/B _5077_/Y _5078_/X vssd1 vssd1 vccd1 vccd1 _5080_/D sky130_fd_sc_hd__o31a_1
XFILLER_29_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8769_ _8769_/A _4361_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[16] sky130_fd_sc_hd__ebufn_8
XFILLER_12_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4450_ _5016_/A vssd1 vssd1 vccd1 vccd1 _4614_/A sky130_fd_sc_hd__clkbuf_2
X_4381_ _4381_/A vssd1 vssd1 vccd1 vccd1 _4381_/Y sky130_fd_sc_hd__inv_2
X_6120_ _5900_/B _5991_/B _5989_/Y vssd1 vssd1 vccd1 vccd1 _6121_/A sky130_fd_sc_hd__a21oi_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6051_ _6169_/A _6051_/B vssd1 vssd1 vccd1 vccd1 _6236_/B sky130_fd_sc_hd__nand2_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5002_ _5117_/A _5147_/B _5002_/C _5002_/D vssd1 vssd1 vccd1 vccd1 _5002_/X sky130_fd_sc_hd__or4_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6953_ _6953_/A _6953_/B vssd1 vssd1 vccd1 vccd1 _6954_/C sky130_fd_sc_hd__xnor2_1
XFILLER_81_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6884_ _6870_/A _6870_/C _6870_/D _6871_/A vssd1 vssd1 vccd1 vccd1 _6884_/X sky130_fd_sc_hd__a22o_1
X_5904_ _6226_/A _5972_/B vssd1 vssd1 vccd1 vccd1 _5905_/B sky130_fd_sc_hd__xor2_1
XFILLER_61_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5835_ _5826_/A _5772_/B _5833_/X _5824_/B vssd1 vssd1 vccd1 vccd1 _5835_/X sky130_fd_sc_hd__a211o_1
XFILLER_34_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8554_ input3/X _8554_/D vssd1 vssd1 vccd1 vccd1 _8554_/Q sky130_fd_sc_hd__dfxtp_1
X_5766_ _5765_/B _5765_/C _5765_/A vssd1 vssd1 vccd1 vccd1 _5776_/B sky130_fd_sc_hd__a21o_1
X_8485_ input3/X _8485_/D vssd1 vssd1 vccd1 vccd1 _8485_/Q sky130_fd_sc_hd__dfxtp_1
X_4717_ _4773_/A vssd1 vssd1 vccd1 vccd1 _4809_/B sky130_fd_sc_hd__clkbuf_2
X_5697_ _5698_/A _5698_/B vssd1 vssd1 vccd1 vccd1 _5812_/B sky130_fd_sc_hd__or2_1
X_7505_ _7505_/A _7505_/B vssd1 vssd1 vccd1 vccd1 _7680_/A sky130_fd_sc_hd__nand2_2
X_4648_ _4711_/A _4649_/B vssd1 vssd1 vccd1 vccd1 _4650_/B sky130_fd_sc_hd__or2_1
X_7436_ _8571_/Q vssd1 vssd1 vccd1 vccd1 _7452_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7367_ _6472_/X _8558_/Q _7362_/X _7366_/X vssd1 vssd1 vccd1 vccd1 _8558_/D sky130_fd_sc_hd__o22a_1
XFILLER_1_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4579_ _6462_/A vssd1 vssd1 vccd1 vccd1 _8410_/A sky130_fd_sc_hd__clkbuf_4
X_6318_ _8536_/Q _8540_/Q _8539_/Q _8535_/Q vssd1 vssd1 vccd1 vccd1 _6320_/B sky130_fd_sc_hd__and4bb_1
X_7298_ _6980_/B _6874_/A _6755_/B _7233_/A vssd1 vssd1 vccd1 vccd1 _7299_/B sky130_fd_sc_hd__o22a_1
XFILLER_1_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6249_ _6249_/A _6249_/B _6249_/C vssd1 vssd1 vccd1 vccd1 _6249_/Y sky130_fd_sc_hd__nand3_1
XFILLER_76_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5620_ _5620_/A _5620_/B _5619_/X vssd1 vssd1 vccd1 vccd1 _5721_/B sky130_fd_sc_hd__or3b_1
X_5551_ _5551_/A _5551_/B vssd1 vssd1 vccd1 vccd1 _5552_/B sky130_fd_sc_hd__nand2_1
X_8270_ _8270_/A _8277_/B vssd1 vssd1 vccd1 vccd1 _8270_/X sky130_fd_sc_hd__or2b_1
X_4502_ _8434_/Q _8433_/Q vssd1 vssd1 vccd1 vccd1 _4516_/A sky130_fd_sc_hd__or2_1
X_7221_ _6914_/A _7038_/A _7206_/B vssd1 vssd1 vccd1 vccd1 _7221_/X sky130_fd_sc_hd__a21o_1
X_5482_ _5493_/A _5497_/B vssd1 vssd1 vccd1 vccd1 _5485_/A sky130_fd_sc_hd__nand2_1
X_4433_ _8464_/Q vssd1 vssd1 vccd1 vccd1 _4761_/B sky130_fd_sc_hd__inv_2
X_4364_ _4382_/A vssd1 vssd1 vccd1 vccd1 _4369_/A sky130_fd_sc_hd__buf_2
X_7152_ _7152_/A _7152_/B vssd1 vssd1 vccd1 vccd1 _7153_/B sky130_fd_sc_hd__nand2_1
X_4295_ _4295_/A vssd1 vssd1 vccd1 vccd1 _4295_/Y sky130_fd_sc_hd__inv_2
X_7083_ _7019_/A _7019_/B _7019_/C _7019_/D vssd1 vssd1 vccd1 vccd1 _7083_/X sky130_fd_sc_hd__a22o_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6103_ _5983_/A _6101_/Y _6102_/Y vssd1 vssd1 vccd1 vccd1 _6114_/A sky130_fd_sc_hd__o21ai_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6034_ _5951_/A _6033_/A _6154_/A vssd1 vssd1 vccd1 vccd1 _6147_/A sky130_fd_sc_hd__a21oi_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7985_ _7982_/B _7983_/Y _7984_/X vssd1 vssd1 vccd1 vccd1 _7986_/B sky130_fd_sc_hd__a21boi_1
XFILLER_26_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6936_ _6904_/Y _6934_/X _6933_/Y _6996_/A vssd1 vssd1 vccd1 vccd1 _6954_/B sky130_fd_sc_hd__o211a_1
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6867_ _7282_/A _6867_/B _6867_/C vssd1 vssd1 vccd1 vccd1 _6871_/A sky130_fd_sc_hd__nand3_1
X_6798_ _7315_/A _6798_/B vssd1 vssd1 vccd1 vccd1 _6891_/A sky130_fd_sc_hd__xor2_1
X_5818_ _5818_/A _5818_/B vssd1 vssd1 vccd1 vccd1 _5818_/Y sky130_fd_sc_hd__nand2_1
XFILLER_22_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8537_ input3/X _8537_/D vssd1 vssd1 vccd1 vccd1 _8537_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5749_ _5746_/B _5749_/B vssd1 vssd1 vccd1 vccd1 _5749_/X sky130_fd_sc_hd__and2b_1
X_8468_ input3/X _8468_/D vssd1 vssd1 vccd1 vccd1 _8468_/Q sky130_fd_sc_hd__dfxtp_4
X_8399_ _8399_/A _8399_/B vssd1 vssd1 vccd1 vccd1 _8401_/A sky130_fd_sc_hd__nor2_1
X_7419_ _8582_/Q vssd1 vssd1 vccd1 vccd1 _8391_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_66_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4982_ _4609_/A _4974_/X _4977_/X _5022_/C _4981_/X vssd1 vssd1 vccd1 vccd1 _4982_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_51_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7770_ _7770_/A _7978_/B vssd1 vssd1 vccd1 vccd1 _8023_/B sky130_fd_sc_hd__nor2_2
X_6721_ _6721_/A _6721_/B vssd1 vssd1 vccd1 vccd1 _6926_/B sky130_fd_sc_hd__xnor2_1
X_6652_ _6652_/A _6652_/B vssd1 vssd1 vccd1 vccd1 _7067_/B sky130_fd_sc_hd__xor2_2
XFILLER_31_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5603_ _5516_/A _5516_/B _5602_/X vssd1 vssd1 vccd1 vccd1 _5635_/A sky130_fd_sc_hd__a21bo_1
X_6583_ _6607_/A vssd1 vssd1 vccd1 vccd1 _6806_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_8322_ _7974_/A _8264_/B _8321_/X vssd1 vssd1 vccd1 vccd1 _8323_/B sky130_fd_sc_hd__a21oi_1
X_5534_ _5649_/A _5543_/A vssd1 vssd1 vccd1 vccd1 _5535_/B sky130_fd_sc_hd__xnor2_2
X_8253_ _8336_/A _8253_/B vssd1 vssd1 vccd1 vccd1 _8255_/C sky130_fd_sc_hd__nand2_1
X_5465_ _5609_/B vssd1 vssd1 vccd1 vccd1 _5518_/C sky130_fd_sc_hd__buf_2
X_7204_ _7180_/A _7180_/B _7180_/C vssd1 vssd1 vccd1 vccd1 _7205_/B sky130_fd_sc_hd__o21ai_1
X_4416_ _5144_/C vssd1 vssd1 vccd1 vccd1 _4466_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_8184_ _8184_/A _8184_/B vssd1 vssd1 vccd1 vccd1 _8186_/B sky130_fd_sc_hd__xor2_1
X_7135_ _7161_/A _7161_/B _7134_/Y vssd1 vssd1 vccd1 vccd1 _7138_/A sky130_fd_sc_hd__a21o_1
X_5396_ _5385_/A _5385_/B _5388_/B _5386_/X vssd1 vssd1 vccd1 vccd1 _5400_/A sky130_fd_sc_hd__a31o_1
X_4347_ _4351_/A vssd1 vssd1 vccd1 vccd1 _4347_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4278_ _4296_/A vssd1 vssd1 vccd1 vccd1 _4283_/A sky130_fd_sc_hd__clkbuf_2
X_7066_ _7122_/C _7148_/B vssd1 vssd1 vccd1 vccd1 _7123_/A sky130_fd_sc_hd__xnor2_1
XTAP_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6017_ _5932_/A _6243_/B _6137_/B vssd1 vssd1 vccd1 vccd1 _6019_/B sky130_fd_sc_hd__a21oi_1
XFILLER_67_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7968_ _8048_/A _8048_/B vssd1 vssd1 vccd1 vccd1 _7976_/A sky130_fd_sc_hd__xor2_2
XFILLER_42_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6919_ _6919_/A _7297_/A vssd1 vssd1 vccd1 vccd1 _6978_/A sky130_fd_sc_hd__xnor2_2
XFILLER_52_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7899_ _7899_/A _8260_/B vssd1 vssd1 vccd1 vccd1 _7899_/X sky130_fd_sc_hd__or2_2
XFILLER_42_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5250_ _8492_/Q _5253_/C vssd1 vssd1 vccd1 vccd1 _5252_/A sky130_fd_sc_hd__and2_1
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5181_ _4623_/X _4642_/A _5179_/Y _5180_/X vssd1 vssd1 vccd1 vccd1 _5181_/X sky130_fd_sc_hd__a31o_1
XFILLER_68_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7822_ _7822_/A _7822_/B vssd1 vssd1 vccd1 vccd1 _8305_/S sky130_fd_sc_hd__nand2_2
X_4965_ _4935_/A _4898_/A _4959_/X _4964_/X vssd1 vssd1 vccd1 vccd1 _4965_/X sky130_fd_sc_hd__o31a_1
X_7753_ _7752_/A _7752_/B _7751_/X vssd1 vssd1 vccd1 vccd1 _7754_/C sky130_fd_sc_hd__o21bai_1
X_6704_ _6705_/A _6705_/B vssd1 vssd1 vccd1 vccd1 _6727_/B sky130_fd_sc_hd__xor2_1
X_4896_ _5064_/A _5153_/A vssd1 vssd1 vccd1 vccd1 _5092_/C sky130_fd_sc_hd__nand2_1
XFILLER_20_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7684_ _7694_/A _7684_/B vssd1 vssd1 vccd1 vccd1 _7702_/A sky130_fd_sc_hd__nand2_1
X_6635_ _7176_/A _7043_/B vssd1 vssd1 vccd1 vccd1 _6919_/A sky130_fd_sc_hd__nor2_1
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6566_ _6647_/A _6784_/A vssd1 vssd1 vccd1 vccd1 _6569_/A sky130_fd_sc_hd__nor2_1
X_5517_ _5601_/B _5517_/B vssd1 vssd1 vccd1 vccd1 _5520_/A sky130_fd_sc_hd__xor2_1
X_8305_ _8306_/A _8123_/A _8305_/S vssd1 vssd1 vccd1 vccd1 _8308_/A sky130_fd_sc_hd__mux2_1
X_6497_ _8552_/Q _8469_/Q vssd1 vssd1 vccd1 vccd1 _6499_/A sky130_fd_sc_hd__and2b_1
X_8236_ _8302_/A _8302_/B vssd1 vssd1 vccd1 vccd1 _8237_/B sky130_fd_sc_hd__xor2_1
X_5448_ _5825_/A vssd1 vssd1 vccd1 vccd1 _5938_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_87_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8167_ _8167_/A _8167_/B vssd1 vssd1 vccd1 vccd1 _8221_/B sky130_fd_sc_hd__xnor2_1
X_5379_ _5417_/A _5404_/B _5378_/X vssd1 vssd1 vccd1 vccd1 _5524_/A sky130_fd_sc_hd__a21o_2
X_7118_ _7118_/A _7118_/B vssd1 vssd1 vccd1 vccd1 _7151_/A sky130_fd_sc_hd__xnor2_2
XFILLER_59_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8098_ _7984_/C _8096_/X _8097_/X vssd1 vssd1 vccd1 vccd1 _8227_/A sky130_fd_sc_hd__o21ai_2
X_7049_ _7106_/A _7106_/B vssd1 vssd1 vccd1 vccd1 _7052_/A sky130_fd_sc_hd__or2b_1
XFILLER_47_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8675__91 vssd1 vssd1 vccd1 vccd1 _8675__91/HI _8784_/A sky130_fd_sc_hd__conb_1
XFILLER_77_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4750_ _4750_/A _4798_/B vssd1 vssd1 vccd1 vccd1 _4885_/A sky130_fd_sc_hd__nor2_2
X_4681_ _4681_/A vssd1 vssd1 vccd1 vccd1 _8467_/D sky130_fd_sc_hd__clkbuf_1
X_6420_ _8554_/Q vssd1 vssd1 vccd1 vccd1 _6455_/A sky130_fd_sc_hd__clkbuf_1
X_6351_ _6351_/A _8534_/Q _6351_/C vssd1 vssd1 vccd1 vccd1 _6357_/C sky130_fd_sc_hd__and3_1
X_5302_ _8507_/Q vssd1 vssd1 vccd1 vccd1 _6281_/B sky130_fd_sc_hd__clkbuf_1
X_6282_ _6282_/A _6282_/B vssd1 vssd1 vccd1 vccd1 _6289_/B sky130_fd_sc_hd__and2_1
X_5233_ _8487_/Q _8486_/Q vssd1 vssd1 vccd1 vccd1 _5234_/C sky130_fd_sc_hd__nand2_1
X_8021_ _7991_/A _7991_/B _7994_/A vssd1 vssd1 vccd1 vccd1 _8086_/A sky130_fd_sc_hd__a21bo_1
X_5164_ _5164_/A _5164_/B _5164_/C _5164_/D vssd1 vssd1 vccd1 vccd1 _5164_/X sky130_fd_sc_hd__or4_1
X_5095_ _5136_/A _5136_/B _5095_/C _5095_/D vssd1 vssd1 vccd1 vccd1 _5095_/X sky130_fd_sc_hd__or4_1
XFILLER_68_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7805_ _7805_/A _7921_/B vssd1 vssd1 vccd1 vccd1 _7808_/A sky130_fd_sc_hd__nand2_2
X_8785_ _8785_/A _4380_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[32] sky130_fd_sc_hd__ebufn_8
XFILLER_52_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5997_ _5984_/A _6183_/S _6002_/A _5804_/B vssd1 vssd1 vccd1 vccd1 _5999_/B sky130_fd_sc_hd__o22a_1
X_4948_ _4935_/X _4942_/X _4947_/X _5112_/B vssd1 vssd1 vccd1 vccd1 _4949_/B sky130_fd_sc_hd__o22ai_1
XFILLER_12_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7736_ _7736_/A _7736_/B _7735_/X vssd1 vssd1 vccd1 vccd1 _7840_/B sky130_fd_sc_hd__or3b_1
X_4879_ _5080_/B _5138_/B vssd1 vssd1 vccd1 vccd1 _4957_/C sky130_fd_sc_hd__or2_1
X_7667_ _7668_/A _7668_/B vssd1 vssd1 vccd1 vccd1 _7715_/A sky130_fd_sc_hd__or2_1
X_6618_ _6804_/B _6618_/B _6618_/C vssd1 vssd1 vccd1 vccd1 _6733_/A sky130_fd_sc_hd__nand3_1
X_7598_ _8317_/A _7969_/A vssd1 vssd1 vccd1 vccd1 _7718_/A sky130_fd_sc_hd__or2_1
X_6549_ _6543_/X _6604_/A _6596_/B _6595_/A _6591_/B vssd1 vssd1 vccd1 vccd1 _6609_/C
+ sky130_fd_sc_hd__a311o_1
XFILLER_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8219_ _8171_/A _8171_/B _8218_/X vssd1 vssd1 vccd1 vccd1 _8295_/A sky130_fd_sc_hd__a21oi_2
XFILLER_87_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5920_ _6006_/A _5921_/B vssd1 vssd1 vccd1 vccd1 _6010_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5851_ _5851_/A _5851_/B vssd1 vssd1 vccd1 vccd1 _5852_/B sky130_fd_sc_hd__nor2_1
X_4802_ _4914_/A _4970_/A vssd1 vssd1 vccd1 vccd1 _5090_/A sky130_fd_sc_hd__or2_2
X_5782_ _5782_/A _5782_/B vssd1 vssd1 vccd1 vccd1 _5783_/B sky130_fd_sc_hd__xor2_4
XFILLER_34_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8570_ input3/X _8570_/D vssd1 vssd1 vccd1 vccd1 _8570_/Q sky130_fd_sc_hd__dfxtp_1
X_4733_ _7506_/B _7501_/B _4737_/A _4738_/B vssd1 vssd1 vccd1 vccd1 _4767_/A sky130_fd_sc_hd__or4_1
X_7521_ _7978_/A vssd1 vssd1 vccd1 vccd1 _7526_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_7452_ _7452_/A _8569_/Q vssd1 vssd1 vccd1 vccd1 _7453_/B sky130_fd_sc_hd__or2b_1
X_6403_ _8563_/Q vssd1 vssd1 vccd1 vccd1 _7384_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_4664_ _4684_/A vssd1 vssd1 vccd1 vccd1 _5192_/B sky130_fd_sc_hd__clkbuf_2
X_4595_ _5121_/B vssd1 vssd1 vccd1 vccd1 _4596_/A sky130_fd_sc_hd__clkbuf_2
X_7383_ _7380_/A _5294_/X _6432_/X _7382_/Y vssd1 vssd1 vccd1 vccd1 _8562_/D sky130_fd_sc_hd__a22o_1
X_6334_ _8528_/Q _8527_/Q _8529_/Q vssd1 vssd1 vccd1 vccd1 _6335_/B sky130_fd_sc_hd__a21o_1
X_6265_ _6251_/X _6264_/X _6261_/X _8519_/Q vssd1 vssd1 vccd1 vccd1 _8519_/D sky130_fd_sc_hd__o2bb2a_1
XFILLER_1_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5216_ _8559_/Q _5202_/A _5215_/X _5213_/X vssd1 vssd1 vccd1 vccd1 _8484_/D sky130_fd_sc_hd__o211a_1
XFILLER_88_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8004_ _8003_/A _8003_/C _8003_/B vssd1 vssd1 vccd1 vccd1 _8005_/B sky130_fd_sc_hd__o21ai_1
X_6196_ _6158_/A _6158_/B _6195_/Y vssd1 vssd1 vccd1 vccd1 _6209_/A sky130_fd_sc_hd__o21a_1
XFILLER_84_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5147_ _5147_/A _5147_/B _5149_/B vssd1 vssd1 vccd1 vccd1 _5147_/X sky130_fd_sc_hd__or3_1
XFILLER_69_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5078_ _4584_/A _5073_/A _4996_/A _5102_/A vssd1 vssd1 vccd1 vccd1 _5078_/X sky130_fd_sc_hd__a211o_1
XFILLER_71_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8768_ _8768_/A _4360_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[15] sky130_fd_sc_hd__ebufn_8
XFILLER_52_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7719_ _7633_/A _7633_/B _7718_/X vssd1 vssd1 vccd1 vccd1 _7754_/A sky130_fd_sc_hd__a21bo_1
XFILLER_40_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8699_ _8699_/A _4279_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[16] sky130_fd_sc_hd__ebufn_8
XFILLER_60_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8645__61 vssd1 vssd1 vccd1 vccd1 _8645__61/HI _8754_/A sky130_fd_sc_hd__conb_1
XFILLER_87_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4380_ _4381_/A vssd1 vssd1 vccd1 vccd1 _4380_/Y sky130_fd_sc_hd__inv_2
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6050_ _6050_/A _5964_/Y vssd1 vssd1 vccd1 vccd1 _6051_/B sky130_fd_sc_hd__or2b_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5001_ _5001_/A _5147_/A vssd1 vssd1 vccd1 vccd1 _5002_/D sky130_fd_sc_hd__or2_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6952_ _6952_/A _6957_/B vssd1 vssd1 vccd1 vccd1 _6953_/B sky130_fd_sc_hd__xnor2_1
XFILLER_53_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6883_ _6883_/A _6883_/B _6883_/C _6883_/D vssd1 vssd1 vccd1 vccd1 _6883_/X sky130_fd_sc_hd__and4_2
X_5903_ _6108_/A _5857_/Y _5902_/X vssd1 vssd1 vccd1 vccd1 _5972_/B sky130_fd_sc_hd__o21a_1
X_5834_ _5823_/Y _5824_/X _5833_/X vssd1 vssd1 vccd1 vccd1 _5836_/A sky130_fd_sc_hd__a21boi_1
XFILLER_34_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8553_ input3/X _8553_/D vssd1 vssd1 vccd1 vccd1 _8553_/Q sky130_fd_sc_hd__dfxtp_1
X_5765_ _5765_/A _5765_/B _5765_/C vssd1 vssd1 vccd1 vccd1 _5776_/A sky130_fd_sc_hd__nand3_1
X_8484_ input3/X _8484_/D vssd1 vssd1 vccd1 vccd1 _8484_/Q sky130_fd_sc_hd__dfxtp_1
X_4716_ _4716_/A vssd1 vssd1 vccd1 vccd1 _4773_/A sky130_fd_sc_hd__clkbuf_2
X_5696_ _5711_/B _5696_/B vssd1 vssd1 vccd1 vccd1 _5698_/B sky130_fd_sc_hd__xnor2_1
X_7504_ _7493_/A _7524_/B _7500_/X _7498_/X vssd1 vssd1 vccd1 vccd1 _7505_/B sky130_fd_sc_hd__a211o_1
X_4647_ _5180_/B vssd1 vssd1 vccd1 vccd1 _4711_/A sky130_fd_sc_hd__clkbuf_2
X_7435_ _7501_/A _8569_/Q vssd1 vssd1 vccd1 vccd1 _7459_/A sky130_fd_sc_hd__and2b_1
X_7366_ _7372_/C _7366_/B _7366_/C vssd1 vssd1 vccd1 vccd1 _7366_/X sky130_fd_sc_hd__and3b_1
XFILLER_89_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6317_ _8530_/Q _8534_/Q _6351_/A _8529_/Q vssd1 vssd1 vccd1 vccd1 _6322_/B sky130_fd_sc_hd__and4bb_1
X_4578_ _7478_/A vssd1 vssd1 vccd1 vccd1 _6462_/A sky130_fd_sc_hd__buf_2
XFILLER_1_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7297_ _7297_/A _7297_/B vssd1 vssd1 vccd1 vccd1 _7299_/A sky130_fd_sc_hd__or2_1
X_6248_ _6248_/A _6254_/B vssd1 vssd1 vccd1 vccd1 _6249_/C sky130_fd_sc_hd__nand2_1
X_6179_ _6179_/A _6162_/A vssd1 vssd1 vccd1 vccd1 _6179_/X sky130_fd_sc_hd__or2b_1
XFILLER_29_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5550_ _5551_/A _5551_/B vssd1 vssd1 vccd1 vccd1 _5599_/A sky130_fd_sc_hd__or2_1
XFILLER_8_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5481_ _8525_/Q _8462_/Q vssd1 vssd1 vccd1 vccd1 _5497_/B sky130_fd_sc_hd__or2b_1
X_4501_ _8440_/Q _8439_/Q _8442_/Q _4501_/D vssd1 vssd1 vccd1 vccd1 _4507_/B sky130_fd_sc_hd__or4_1
X_7220_ _7183_/A _7121_/A _7184_/C _7248_/A vssd1 vssd1 vccd1 vccd1 _7232_/A sky130_fd_sc_hd__o22a_1
X_4432_ _4762_/A vssd1 vssd1 vccd1 vccd1 _4759_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7151_ _7151_/A _7151_/B vssd1 vssd1 vccd1 vccd1 _7193_/B sky130_fd_sc_hd__xor2_2
X_4363_ _4363_/A vssd1 vssd1 vccd1 vccd1 _4363_/Y sky130_fd_sc_hd__inv_2
X_4294_ _4295_/A vssd1 vssd1 vccd1 vccd1 _4294_/Y sky130_fd_sc_hd__inv_2
X_7082_ _7136_/A _7136_/B vssd1 vssd1 vccd1 vccd1 _7082_/X sky130_fd_sc_hd__and2_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6102_ _6104_/A _6102_/B vssd1 vssd1 vccd1 vccd1 _6102_/Y sky130_fd_sc_hd__nand2_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6033_ _6033_/A _6153_/C vssd1 vssd1 vccd1 vccd1 _6154_/B sky130_fd_sc_hd__xnor2_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7984_ _7984_/A _8105_/A _7984_/C vssd1 vssd1 vccd1 vccd1 _7984_/X sky130_fd_sc_hd__or3_1
XFILLER_81_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6935_ _6996_/A _6933_/Y _6934_/X _6904_/Y vssd1 vssd1 vccd1 vccd1 _6954_/A sky130_fd_sc_hd__a211oi_4
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6866_ _6848_/A _6848_/B _6848_/C vssd1 vssd1 vccd1 vccd1 _6867_/C sky130_fd_sc_hd__a21o_1
XFILLER_34_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6797_ _7310_/S _6708_/B _6796_/Y vssd1 vssd1 vccd1 vccd1 _6798_/B sky130_fd_sc_hd__a21o_1
XFILLER_10_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5817_ _6061_/A _6061_/B _5816_/X vssd1 vssd1 vccd1 vccd1 _5893_/A sky130_fd_sc_hd__a21o_1
X_8536_ input3/X _8536_/D vssd1 vssd1 vccd1 vccd1 _8536_/Q sky130_fd_sc_hd__dfxtp_1
X_5748_ _5892_/A _5748_/B vssd1 vssd1 vccd1 vccd1 _6057_/B sky130_fd_sc_hd__xnor2_1
XFILLER_22_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8467_ input3/X _8467_/D vssd1 vssd1 vccd1 vccd1 _8467_/Q sky130_fd_sc_hd__dfxtp_2
X_5679_ _5577_/A _5679_/B vssd1 vssd1 vccd1 vccd1 _6090_/D sky130_fd_sc_hd__and2b_1
X_7418_ _8583_/Q vssd1 vssd1 vccd1 vccd1 _8397_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_8398_ _8397_/B _8412_/B vssd1 vssd1 vccd1 vccd1 _8399_/B sky130_fd_sc_hd__and2b_1
X_7349_ _7349_/A _7349_/B vssd1 vssd1 vccd1 vccd1 _7372_/A sky130_fd_sc_hd__xor2_2
XFILLER_1_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8615__31 vssd1 vssd1 vccd1 vccd1 _8615__31/HI _8710_/A sky130_fd_sc_hd__conb_1
XFILLER_66_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4981_ _5016_/A _5112_/D _4981_/C vssd1 vssd1 vccd1 vccd1 _4981_/X sky130_fd_sc_hd__or3_1
X_6720_ _6700_/B _6700_/C _6700_/A vssd1 vssd1 vccd1 vccd1 _6725_/C sky130_fd_sc_hd__a21oi_1
X_6651_ _6939_/B _6714_/C _6672_/A vssd1 vssd1 vccd1 vccd1 _6657_/A sky130_fd_sc_hd__or3_4
X_6582_ _6660_/A _6929_/B vssd1 vssd1 vccd1 vccd1 _6930_/A sky130_fd_sc_hd__nand2_1
X_5602_ _5602_/A _5505_/B vssd1 vssd1 vccd1 vccd1 _5602_/X sky130_fd_sc_hd__or2b_1
X_8321_ _8263_/A _8321_/B vssd1 vssd1 vccd1 vccd1 _8321_/X sky130_fd_sc_hd__and2b_1
X_5533_ _5648_/A _5984_/A vssd1 vssd1 vccd1 vccd1 _5543_/A sky130_fd_sc_hd__nor2_2
X_8252_ _8252_/A _8252_/B vssd1 vssd1 vccd1 vccd1 _8253_/B sky130_fd_sc_hd__or2_1
X_5464_ _5492_/B _5467_/A vssd1 vssd1 vccd1 vccd1 _5609_/B sky130_fd_sc_hd__or2_1
X_7203_ _6714_/A _7185_/A _7202_/Y _7070_/B vssd1 vssd1 vccd1 vccd1 _7219_/A sky130_fd_sc_hd__o22a_1
X_4415_ _7506_/B vssd1 vssd1 vccd1 vccd1 _5144_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_5395_ _5685_/A _6244_/B vssd1 vssd1 vccd1 vccd1 _5410_/A sky130_fd_sc_hd__nand2_1
X_8183_ _8194_/A _8194_/B _8182_/X vssd1 vssd1 vccd1 vccd1 _8186_/A sky130_fd_sc_hd__a21oi_1
X_4346_ _4358_/A vssd1 vssd1 vccd1 vccd1 _4351_/A sky130_fd_sc_hd__buf_2
X_7134_ _7134_/A _7134_/B vssd1 vssd1 vccd1 vccd1 _7134_/Y sky130_fd_sc_hd__nor2_1
XFILLER_86_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4277_ _4277_/A vssd1 vssd1 vccd1 vccd1 _4277_/Y sky130_fd_sc_hd__inv_2
X_7065_ _7065_/A _7065_/B vssd1 vssd1 vccd1 vccd1 _7136_/A sky130_fd_sc_hd__nor2_1
XFILLER_86_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6016_ _5945_/A _6014_/X _6015_/X vssd1 vssd1 vccd1 vccd1 _6124_/A sky130_fd_sc_hd__a21oi_2
XFILLER_36_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7967_ _7967_/A _7967_/B vssd1 vssd1 vccd1 vccd1 _8048_/B sky130_fd_sc_hd__xnor2_1
XFILLER_42_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6918_ _6918_/A _6917_/X vssd1 vssd1 vccd1 vccd1 _6921_/A sky130_fd_sc_hd__or2b_1
X_7898_ _7898_/A _7898_/B vssd1 vssd1 vccd1 vccd1 _7944_/A sky130_fd_sc_hd__and2_2
X_6849_ _6914_/C _6554_/Y vssd1 vssd1 vccd1 vccd1 _6850_/A sky130_fd_sc_hd__or2b_1
XFILLER_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8519_ input3/X _8519_/D vssd1 vssd1 vccd1 vccd1 _8519_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5180_ _5180_/A _5180_/B _4655_/A vssd1 vssd1 vccd1 vccd1 _5180_/X sky130_fd_sc_hd__or3b_1
XFILLER_95_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7821_ _8176_/A _8176_/B vssd1 vssd1 vccd1 vccd1 _7834_/A sky130_fd_sc_hd__and2_1
X_4964_ _5135_/A _4906_/B _4939_/B _4962_/X _4963_/X vssd1 vssd1 vccd1 vccd1 _4964_/X
+ sky130_fd_sc_hd__a2111o_1
X_7752_ _7752_/A _7752_/B _7751_/X vssd1 vssd1 vccd1 vccd1 _7839_/B sky130_fd_sc_hd__or3b_1
X_6703_ _6703_/A _6703_/B vssd1 vssd1 vccd1 vccd1 _6705_/B sky130_fd_sc_hd__xor2_1
XFILLER_51_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4895_ _5093_/A vssd1 vssd1 vccd1 vccd1 _5153_/A sky130_fd_sc_hd__clkbuf_2
X_7683_ _8367_/A _7530_/A _8101_/C _7682_/Y _7533_/X vssd1 vssd1 vccd1 vccd1 _7684_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_32_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6634_ _6751_/A vssd1 vssd1 vccd1 vccd1 _7176_/A sky130_fd_sc_hd__clkbuf_2
X_6565_ _6693_/C vssd1 vssd1 vccd1 vccd1 _6784_/A sky130_fd_sc_hd__clkbuf_2
X_6496_ _6501_/A _6501_/B _6495_/X vssd1 vssd1 vccd1 vccd1 _6500_/A sky130_fd_sc_hd__a21o_2
X_8304_ _8235_/A _8235_/B _8234_/A vssd1 vssd1 vccd1 vccd1 _8309_/A sky130_fd_sc_hd__a21oi_1
X_5516_ _5516_/A _5516_/B vssd1 vssd1 vccd1 vccd1 _5517_/B sky130_fd_sc_hd__xnor2_1
X_8235_ _8235_/A _8235_/B vssd1 vssd1 vccd1 vccd1 _8302_/B sky130_fd_sc_hd__xor2_1
X_5447_ _5615_/A vssd1 vssd1 vccd1 vccd1 _5825_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_59_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8166_ _8166_/A _8166_/B vssd1 vssd1 vccd1 vccd1 _8167_/B sky130_fd_sc_hd__nor2_1
X_5378_ _8510_/Q _7498_/B vssd1 vssd1 vccd1 vccd1 _5378_/X sky130_fd_sc_hd__and2b_1
X_4329_ _4332_/A vssd1 vssd1 vccd1 vccd1 _4329_/Y sky130_fd_sc_hd__inv_2
X_7117_ _7250_/A _6657_/A _7116_/Y vssd1 vssd1 vccd1 vccd1 _7118_/B sky130_fd_sc_hd__o21a_1
X_8097_ _8097_/A _8249_/B vssd1 vssd1 vccd1 vccd1 _8097_/X sky130_fd_sc_hd__or2_1
X_7048_ _7057_/A _7057_/B vssd1 vssd1 vccd1 vccd1 _7106_/B sky130_fd_sc_hd__xor2_1
XFILLER_59_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4680_ _8403_/A _4680_/B vssd1 vssd1 vccd1 vccd1 _4681_/A sky130_fd_sc_hd__and2_1
X_6350_ _6350_/A _6350_/B vssd1 vssd1 vccd1 vccd1 _8533_/D sky130_fd_sc_hd__nor2_1
X_5301_ _8523_/Q vssd1 vssd1 vccd1 vccd1 _6281_/A sky130_fd_sc_hd__inv_2
X_6281_ _6281_/A _6281_/B vssd1 vssd1 vccd1 vccd1 _6282_/B sky130_fd_sc_hd__or2_1
X_5232_ _5260_/A vssd1 vssd1 vccd1 vccd1 _5291_/A sky130_fd_sc_hd__clkbuf_2
X_8020_ _8013_/A _8013_/B _8019_/X vssd1 vssd1 vccd1 vccd1 _8084_/A sky130_fd_sc_hd__a21oi_1
X_5163_ _4973_/A _5148_/A _5169_/D _5156_/A vssd1 vssd1 vccd1 vccd1 _5164_/D sky130_fd_sc_hd__a211o_1
XFILLER_68_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5094_ _5019_/A _5117_/A _5022_/B _5093_/X vssd1 vssd1 vccd1 vccd1 _5095_/D sky130_fd_sc_hd__o31a_1
XFILLER_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7804_ _7804_/A _7983_/B _7804_/C vssd1 vssd1 vccd1 vccd1 _7810_/B sky130_fd_sc_hd__and3_1
XFILLER_37_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8784_ _8784_/A _4379_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[31] sky130_fd_sc_hd__ebufn_8
X_5996_ _5957_/A _5957_/B _5995_/X vssd1 vssd1 vccd1 vccd1 _6098_/A sky130_fd_sc_hd__a21oi_1
X_4947_ _5146_/A _4987_/A _4947_/C _4947_/D vssd1 vssd1 vccd1 vccd1 _4947_/X sky130_fd_sc_hd__or4_1
XFILLER_52_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7735_ _7860_/A _7860_/B vssd1 vssd1 vccd1 vccd1 _7735_/X sky130_fd_sc_hd__xor2_1
X_4878_ _5010_/A vssd1 vssd1 vccd1 vccd1 _5171_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7666_ _7654_/B _7547_/Y _7656_/B vssd1 vssd1 vccd1 vccd1 _7668_/B sky130_fd_sc_hd__o21ai_1
X_6617_ _6616_/B _6616_/C _6804_/A vssd1 vssd1 vccd1 vccd1 _6618_/C sky130_fd_sc_hd__a21o_1
X_7597_ _7962_/A vssd1 vssd1 vccd1 vccd1 _8317_/A sky130_fd_sc_hd__clkbuf_2
X_6548_ _8555_/Q _7539_/B vssd1 vssd1 vccd1 vccd1 _6591_/B sky130_fd_sc_hd__nor2_1
XFILLER_3_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6479_ _6479_/A _6479_/B vssd1 vssd1 vccd1 vccd1 _6999_/B sky130_fd_sc_hd__nor2_2
X_8218_ _8170_/B _8218_/B vssd1 vssd1 vccd1 vccd1 _8218_/X sky130_fd_sc_hd__and2b_1
XFILLER_87_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_0 _7185_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8149_ _8260_/C _8149_/B vssd1 vssd1 vccd1 vccd1 _8258_/B sky130_fd_sc_hd__xnor2_1
XFILLER_75_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5850_ _5851_/A _5851_/B vssd1 vssd1 vccd1 vccd1 _5923_/A sky130_fd_sc_hd__and2_2
XFILLER_34_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4801_ _5020_/B _4915_/A vssd1 vssd1 vccd1 vccd1 _4970_/A sky130_fd_sc_hd__or2_1
XFILLER_61_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5781_ _5781_/A _5781_/B vssd1 vssd1 vccd1 vccd1 _5782_/B sky130_fd_sc_hd__xnor2_4
X_4732_ _4976_/A _4975_/B vssd1 vssd1 vccd1 vccd1 _5138_/A sky130_fd_sc_hd__or2_2
XFILLER_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7520_ _7520_/A _7520_/B vssd1 vssd1 vccd1 vccd1 _7978_/A sky130_fd_sc_hd__xnor2_4
X_4663_ _4663_/A _4663_/B vssd1 vssd1 vccd1 vccd1 _4684_/A sky130_fd_sc_hd__and2_1
XFILLER_9_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7451_ _8569_/Q _7452_/A vssd1 vssd1 vccd1 vccd1 _7453_/A sky130_fd_sc_hd__or2b_1
X_6402_ _7410_/A _6424_/B _7403_/B vssd1 vssd1 vccd1 vccd1 _6402_/Y sky130_fd_sc_hd__o21ai_1
X_4594_ _5064_/A _4945_/A vssd1 vssd1 vccd1 vccd1 _5121_/B sky130_fd_sc_hd__nand2_1
X_7382_ _8561_/Q _7382_/B vssd1 vssd1 vccd1 vccd1 _7382_/Y sky130_fd_sc_hd__xnor2_1
X_6333_ _8529_/Q _8528_/Q _8527_/Q vssd1 vssd1 vccd1 vccd1 _6338_/B sky130_fd_sc_hd__and3_1
XFILLER_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6264_ _6264_/A _6264_/B _6264_/C _6264_/D vssd1 vssd1 vccd1 vccd1 _6264_/X sky130_fd_sc_hd__or4_1
X_5215_ _8484_/Q _5217_/B vssd1 vssd1 vccd1 vccd1 _5215_/X sky130_fd_sc_hd__or2_1
X_8003_ _8003_/A _8003_/B _8003_/C vssd1 vssd1 vccd1 vccd1 _8003_/Y sky130_fd_sc_hd__nor3_1
X_6195_ _6195_/A _6195_/B vssd1 vssd1 vccd1 vccd1 _6195_/Y sky130_fd_sc_hd__nand2_1
XFILLER_84_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5146_ _5146_/A _5149_/B _5146_/C _5160_/D vssd1 vssd1 vccd1 vccd1 _5146_/X sky130_fd_sc_hd__or4_1
XFILLER_56_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5077_ _4584_/A _4791_/A _5088_/A vssd1 vssd1 vccd1 vccd1 _5077_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_84_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8767_ _8767_/A _4359_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[14] sky130_fd_sc_hd__ebufn_8
XFILLER_52_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5979_ _5980_/C _6106_/A _5579_/B vssd1 vssd1 vccd1 vccd1 _5981_/B sky130_fd_sc_hd__a21o_1
X_7718_ _7718_/A _7624_/B vssd1 vssd1 vccd1 vccd1 _7718_/X sky130_fd_sc_hd__or2b_1
XFILLER_40_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8698_ _8698_/A _4277_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[15] sky130_fd_sc_hd__ebufn_8
X_7649_ _7649_/A _7649_/B vssd1 vssd1 vccd1 vccd1 _8105_/A sky130_fd_sc_hd__xnor2_4
XFILLER_4_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8660__76 vssd1 vssd1 vccd1 vccd1 _8660__76/HI _8769_/A sky130_fd_sc_hd__conb_1
XFILLER_47_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5000_ _4955_/A _4938_/A _5089_/B _4945_/Y _4898_/A vssd1 vssd1 vccd1 vccd1 _5002_/C
+ sky130_fd_sc_hd__o32a_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6951_ _7310_/S _6951_/B vssd1 vssd1 vccd1 vccd1 _6957_/B sky130_fd_sc_hd__xnor2_1
XFILLER_81_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6882_ _6880_/A _6880_/C _6880_/B vssd1 vssd1 vccd1 vccd1 _6883_/D sky130_fd_sc_hd__a21o_1
X_5902_ _5902_/A _6126_/B vssd1 vssd1 vccd1 vccd1 _5902_/X sky130_fd_sc_hd__or2_1
XFILLER_46_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5833_ _5833_/A _5833_/B vssd1 vssd1 vccd1 vccd1 _5833_/X sky130_fd_sc_hd__xor2_1
XFILLER_34_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8552_ input3/X _8552_/D vssd1 vssd1 vccd1 vccd1 _8552_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5764_ _5764_/A _5764_/B _5764_/C _5943_/A vssd1 vssd1 vccd1 vccd1 _5765_/C sky130_fd_sc_hd__or4_2
X_7503_ _7641_/A _7641_/B vssd1 vssd1 vccd1 vccd1 _7805_/A sky130_fd_sc_hd__xor2_4
X_8483_ input3/X _8483_/D vssd1 vssd1 vccd1 vccd1 _8483_/Q sky130_fd_sc_hd__dfxtp_1
X_4715_ _4715_/A _4737_/A _4738_/B _5144_/C vssd1 vssd1 vccd1 vccd1 _4716_/A sky130_fd_sc_hd__or4b_1
X_5695_ _5805_/A _5860_/A vssd1 vssd1 vccd1 vccd1 _5696_/B sky130_fd_sc_hd__nor2_1
X_4646_ _4646_/A vssd1 vssd1 vccd1 vccd1 _8460_/D sky130_fd_sc_hd__clkbuf_1
X_7434_ _8572_/Q vssd1 vssd1 vccd1 vccd1 _7501_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7365_ _7365_/A _7365_/B vssd1 vssd1 vccd1 vccd1 _7366_/C sky130_fd_sc_hd__nand2_1
X_4577_ _6427_/A vssd1 vssd1 vccd1 vccd1 _7478_/A sky130_fd_sc_hd__buf_4
X_6316_ _8528_/Q _8527_/Q vssd1 vssd1 vccd1 vccd1 _6322_/A sky130_fd_sc_hd__nor2_1
XFILLER_89_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7296_ _7296_/A _7296_/B vssd1 vssd1 vccd1 vccd1 _7300_/A sky130_fd_sc_hd__or2_1
XFILLER_1_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6247_ _6247_/A _6247_/B vssd1 vssd1 vccd1 vccd1 _6254_/B sky130_fd_sc_hd__xnor2_1
XFILLER_57_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6178_ _6162_/A _6179_/A vssd1 vssd1 vccd1 vccd1 _6178_/X sky130_fd_sc_hd__and2b_1
X_5129_ _5178_/B _4639_/A _4711_/B vssd1 vssd1 vccd1 vccd1 _5130_/S sky130_fd_sc_hd__o21a_1
XFILLER_72_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4500_ _8444_/Q _8443_/Q _8446_/Q _8445_/Q vssd1 vssd1 vccd1 vccd1 _4501_/D sky130_fd_sc_hd__or4_1
XFILLER_8_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5480_ _6514_/A _6293_/A vssd1 vssd1 vccd1 vccd1 _5493_/A sky130_fd_sc_hd__or2b_1
X_4431_ _8465_/Q vssd1 vssd1 vccd1 vccd1 _4762_/A sky130_fd_sc_hd__inv_2
XFILLER_6_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7150_ _7181_/A _7181_/B vssd1 vssd1 vccd1 vccd1 _7193_/A sky130_fd_sc_hd__and2_1
X_4362_ _4363_/A vssd1 vssd1 vccd1 vccd1 _4362_/Y sky130_fd_sc_hd__inv_2
X_4293_ _4295_/A vssd1 vssd1 vccd1 vccd1 _4293_/Y sky130_fd_sc_hd__inv_2
X_7081_ _7081_/A _7081_/B vssd1 vssd1 vccd1 vccd1 _7136_/B sky130_fd_sc_hd__xor2_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6101_ _6101_/A vssd1 vssd1 vccd1 vccd1 _6101_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6032_ _6151_/S _6032_/B vssd1 vssd1 vccd1 vccd1 _6153_/C sky130_fd_sc_hd__xnor2_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7983_ _7983_/A _7983_/B vssd1 vssd1 vccd1 vccd1 _7983_/Y sky130_fd_sc_hd__nand2_1
X_6934_ _6904_/A _6904_/C _6904_/B vssd1 vssd1 vccd1 vccd1 _6934_/X sky130_fd_sc_hd__o21a_1
XFILLER_54_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6865_ _6874_/A _6874_/B _6874_/C vssd1 vssd1 vccd1 vccd1 _6867_/B sky130_fd_sc_hd__and3_1
XFILLER_34_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6796_ _6796_/A _6796_/B vssd1 vssd1 vccd1 vccd1 _6796_/Y sky130_fd_sc_hd__nor2_1
XFILLER_10_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5816_ _5815_/B _5816_/B vssd1 vssd1 vccd1 vccd1 _5816_/X sky130_fd_sc_hd__and2b_1
X_8535_ input3/X _8535_/D vssd1 vssd1 vccd1 vccd1 _8535_/Q sky130_fd_sc_hd__dfxtp_1
X_5747_ _5812_/B _5747_/B vssd1 vssd1 vccd1 vccd1 _5892_/A sky130_fd_sc_hd__nand2_1
XFILLER_10_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8589__5 vssd1 vssd1 vccd1 vccd1 _8589__5/HI _8684_/A sky130_fd_sc_hd__conb_1
X_8466_ input3/X _8466_/D vssd1 vssd1 vccd1 vccd1 _8466_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5678_ _6087_/A _6090_/B vssd1 vssd1 vccd1 vccd1 _6083_/B sky130_fd_sc_hd__nor2b_1
X_7417_ _7417_/A vssd1 vssd1 vccd1 vccd1 _7417_/Y sky130_fd_sc_hd__inv_2
X_4629_ _4629_/A _5175_/S vssd1 vssd1 vccd1 vccd1 _4629_/Y sky130_fd_sc_hd__nand2_1
X_8397_ _8412_/B _8397_/B vssd1 vssd1 vccd1 vccd1 _8399_/A sky130_fd_sc_hd__and2b_1
X_7348_ _7338_/X _7339_/Y _7342_/Y _7344_/X _7347_/Y vssd1 vssd1 vccd1 vccd1 _7356_/C
+ sky130_fd_sc_hd__o2111a_1
X_7279_ _7279_/A _7279_/B vssd1 vssd1 vccd1 vccd1 _7335_/A sky130_fd_sc_hd__xnor2_1
XFILLER_1_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8630__46 vssd1 vssd1 vccd1 vccd1 _8630__46/HI _8725_/A sky130_fd_sc_hd__conb_1
XFILLER_82_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4980_ _5112_/A _4941_/D _5022_/B _5089_/B _4920_/X vssd1 vssd1 vccd1 vccd1 _4981_/C
+ sky130_fd_sc_hd__o32a_1
XFILLER_51_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6650_ _6682_/A _6682_/B vssd1 vssd1 vccd1 vccd1 _6672_/A sky130_fd_sc_hd__xnor2_2
XFILLER_31_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6581_ _6702_/A _6581_/B vssd1 vssd1 vccd1 vccd1 _6929_/B sky130_fd_sc_hd__xnor2_1
X_5601_ _5517_/B _5601_/B vssd1 vssd1 vccd1 vccd1 _5639_/A sky130_fd_sc_hd__and2b_1
X_8320_ _8278_/A _8279_/A _8278_/B vssd1 vssd1 vccd1 vccd1 _8324_/A sky130_fd_sc_hd__o21ba_1
X_5532_ _5532_/A _5532_/B vssd1 vssd1 vccd1 vccd1 _5984_/A sky130_fd_sc_hd__xnor2_4
XFILLER_8_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8251_ _8252_/A _8252_/B vssd1 vssd1 vccd1 vccd1 _8336_/A sky130_fd_sc_hd__nand2_1
X_5463_ _5463_/A _5463_/B vssd1 vssd1 vccd1 vccd1 _5467_/A sky130_fd_sc_hd__xnor2_1
X_5394_ _5648_/A vssd1 vssd1 vccd1 vccd1 _6244_/B sky130_fd_sc_hd__clkbuf_2
X_8182_ _8181_/A _8182_/B vssd1 vssd1 vccd1 vccd1 _8182_/X sky130_fd_sc_hd__and2b_1
X_7202_ _7202_/A _7202_/B vssd1 vssd1 vccd1 vccd1 _7202_/Y sky130_fd_sc_hd__nor2_1
X_4414_ _8470_/Q vssd1 vssd1 vccd1 vccd1 _7506_/B sky130_fd_sc_hd__clkbuf_4
X_7133_ _7133_/A _7133_/B vssd1 vssd1 vccd1 vccd1 _7161_/B sky130_fd_sc_hd__xor2_1
X_4345_ _4345_/A vssd1 vssd1 vccd1 vccd1 _4345_/Y sky130_fd_sc_hd__inv_2
X_7064_ _7064_/A _7064_/B _7064_/C vssd1 vssd1 vccd1 vccd1 _7065_/B sky130_fd_sc_hd__and3_1
X_4276_ _4277_/A vssd1 vssd1 vccd1 vccd1 _4276_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6015_ _6015_/A _6015_/B vssd1 vssd1 vccd1 vccd1 _6015_/X sky130_fd_sc_hd__and2_1
XFILLER_39_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7966_ _7966_/A _7966_/B vssd1 vssd1 vccd1 vccd1 _7967_/B sky130_fd_sc_hd__xor2_2
X_6917_ _6916_/A _6916_/C _6916_/B vssd1 vssd1 vccd1 vccd1 _6917_/X sky130_fd_sc_hd__a21o_1
XFILLER_54_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7897_ _7861_/A _7888_/X _7862_/B _7896_/Y vssd1 vssd1 vccd1 vccd1 _7902_/A sky130_fd_sc_hd__a2bb2o_2
XFILLER_23_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6848_ _6848_/A _6848_/B _6848_/C vssd1 vssd1 vccd1 vccd1 _7282_/A sky130_fd_sc_hd__nand3_2
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6779_ _6764_/A _6764_/B _6778_/Y vssd1 vssd1 vccd1 vccd1 _6783_/A sky130_fd_sc_hd__o21a_1
X_8518_ input3/X _8518_/D vssd1 vssd1 vccd1 vccd1 _8518_/Q sky130_fd_sc_hd__dfxtp_1
X_8449_ input3/X _8449_/D vssd1 vssd1 vccd1 vccd1 _8449_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7820_ _7933_/B _7871_/B _7872_/B vssd1 vssd1 vccd1 vccd1 _7836_/A sky130_fd_sc_hd__and3_1
XFILLER_36_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4963_ _4848_/A _4885_/A _5088_/A vssd1 vssd1 vccd1 vccd1 _4963_/X sky130_fd_sc_hd__a21o_1
X_7751_ _7838_/A _7751_/B vssd1 vssd1 vccd1 vccd1 _7751_/X sky130_fd_sc_hd__and2_1
X_6702_ _6702_/A _6581_/B vssd1 vssd1 vccd1 vccd1 _6705_/A sky130_fd_sc_hd__or2b_1
XFILLER_51_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7682_ _7682_/A _7682_/B vssd1 vssd1 vccd1 vccd1 _7682_/Y sky130_fd_sc_hd__nand2_1
X_4894_ _5089_/A vssd1 vssd1 vccd1 vccd1 _5135_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6633_ _6626_/Y _6755_/A vssd1 vssd1 vccd1 vccd1 _6892_/A sky130_fd_sc_hd__and2b_1
XFILLER_32_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6564_ _6652_/A _6652_/B vssd1 vssd1 vccd1 vccd1 _6693_/C sky130_fd_sc_hd__xnor2_1
X_6495_ _8551_/Q _8468_/Q vssd1 vssd1 vccd1 vccd1 _6495_/X sky130_fd_sc_hd__and2b_1
X_8303_ _8237_/A _8237_/B _8302_/Y vssd1 vssd1 vccd1 vccd1 _8310_/A sky130_fd_sc_hd__a21bo_1
X_5515_ _5778_/A _5637_/B _5515_/C vssd1 vssd1 vccd1 vccd1 _5516_/B sky130_fd_sc_hd__and3b_1
X_8234_ _8234_/A _8234_/B vssd1 vssd1 vccd1 vccd1 _8235_/B sky130_fd_sc_hd__nor2_1
X_5446_ _5609_/A vssd1 vssd1 vccd1 vccd1 _5615_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_87_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8165_ _8165_/A _8165_/B _8165_/C vssd1 vssd1 vccd1 vccd1 _8166_/B sky130_fd_sc_hd__nor3_1
X_5377_ _8510_/Q _8468_/Q vssd1 vssd1 vccd1 vccd1 _5404_/B sky130_fd_sc_hd__xnor2_4
X_4328_ _4332_/A vssd1 vssd1 vccd1 vccd1 _4328_/Y sky130_fd_sc_hd__inv_2
X_8096_ _8097_/A _8249_/B vssd1 vssd1 vccd1 vccd1 _8096_/X sky130_fd_sc_hd__and2_1
X_7116_ _7116_/A _7116_/B vssd1 vssd1 vccd1 vccd1 _7116_/Y sky130_fd_sc_hd__nand2_1
X_7047_ _7099_/B _7099_/C _7099_/A vssd1 vssd1 vccd1 vccd1 _7057_/B sky130_fd_sc_hd__a21bo_1
XFILLER_59_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4259_ _4390_/A vssd1 vssd1 vccd1 vccd1 _4264_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_27_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8600__16 vssd1 vssd1 vccd1 vccd1 _8600__16/HI _8695_/A sky130_fd_sc_hd__conb_1
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7949_ _8326_/A _7949_/B vssd1 vssd1 vccd1 vccd1 _7956_/A sky130_fd_sc_hd__xnor2_1
XFILLER_27_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5300_ _6274_/B _6270_/A _8523_/Q vssd1 vssd1 vccd1 vccd1 _5300_/X sky130_fd_sc_hd__o21a_1
X_6280_ _6276_/B _6278_/B _6276_/A vssd1 vssd1 vccd1 vccd1 _6282_/A sky130_fd_sc_hd__o21ba_1
XFILLER_69_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5231_ _5231_/A vssd1 vssd1 vccd1 vccd1 _8486_/D sky130_fd_sc_hd__clkbuf_1
X_8666__82 vssd1 vssd1 vccd1 vccd1 _8666__82/HI _8775_/A sky130_fd_sc_hd__conb_1
X_5162_ _5162_/A _5162_/B vssd1 vssd1 vccd1 vccd1 _5169_/D sky130_fd_sc_hd__or2_1
X_5093_ _5093_/A _5093_/B _5093_/C _5093_/D vssd1 vssd1 vccd1 vccd1 _5093_/X sky130_fd_sc_hd__or4_1
XFILLER_96_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8783_ _8783_/A _4378_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[30] sky130_fd_sc_hd__ebufn_8
X_7803_ _7803_/A vssd1 vssd1 vccd1 vccd1 _7983_/B sky130_fd_sc_hd__clkbuf_2
X_5995_ _5956_/A _5995_/B vssd1 vssd1 vccd1 vccd1 _5995_/X sky130_fd_sc_hd__and2b_1
X_7734_ _7734_/A _7746_/A vssd1 vssd1 vccd1 vccd1 _7860_/B sky130_fd_sc_hd__xnor2_1
X_4946_ _4839_/A _5151_/B _5164_/A _4945_/Y _4989_/A vssd1 vssd1 vccd1 vccd1 _4947_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_33_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4877_ _5102_/A vssd1 vssd1 vccd1 vccd1 _5088_/A sky130_fd_sc_hd__buf_2
X_7665_ _7665_/A _7665_/B vssd1 vssd1 vccd1 vccd1 _7668_/A sky130_fd_sc_hd__nand2_1
X_6616_ _6804_/A _6616_/B _6616_/C vssd1 vssd1 vccd1 vccd1 _6618_/B sky130_fd_sc_hd__nand3_1
X_7596_ _7731_/A vssd1 vssd1 vccd1 vccd1 _7962_/A sky130_fd_sc_hd__clkbuf_1
X_6547_ _8554_/Q _8471_/Q vssd1 vssd1 vccd1 vccd1 _6595_/A sky130_fd_sc_hd__and2b_1
XFILLER_20_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6478_ _8459_/Q _8563_/Q vssd1 vssd1 vccd1 vccd1 _6479_/B sky130_fd_sc_hd__and2b_1
X_8217_ _8192_/X _8355_/A _8355_/B _8216_/X vssd1 vssd1 vccd1 vccd1 _8364_/B sky130_fd_sc_hd__a31o_1
X_5429_ _5429_/A _5429_/B vssd1 vssd1 vccd1 vccd1 _5560_/A sky130_fd_sc_hd__xnor2_1
XFILLER_87_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8148_ _8148_/A _8154_/A vssd1 vssd1 vccd1 vccd1 _8149_/B sky130_fd_sc_hd__xor2_2
XINSDIODE2_1 _7194_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8079_ _8088_/A _8088_/B vssd1 vssd1 vccd1 vccd1 _8080_/B sky130_fd_sc_hd__xor2_1
XFILLER_74_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4800_ _4800_/A _4953_/B vssd1 vssd1 vccd1 vccd1 _4915_/A sky130_fd_sc_hd__nor2_1
XFILLER_21_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5780_ _5823_/A _5780_/B vssd1 vssd1 vccd1 vccd1 _5781_/B sky130_fd_sc_hd__xor2_4
XFILLER_34_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4731_ _4809_/B _4782_/B _5169_/A vssd1 vssd1 vccd1 vccd1 _4975_/B sky130_fd_sc_hd__o21bai_2
XFILLER_14_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4662_ _4754_/B _4663_/B _4661_/X vssd1 vssd1 vccd1 vccd1 _8464_/D sky130_fd_sc_hd__a21oi_1
X_7450_ _7494_/A _7448_/X _7449_/Y vssd1 vssd1 vccd1 vccd1 _8570_/D sky130_fd_sc_hd__o21a_1
X_6401_ _7390_/A vssd1 vssd1 vccd1 vccd1 _7403_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_4593_ _4593_/A _6521_/B _5441_/B vssd1 vssd1 vccd1 vccd1 _4659_/B sky130_fd_sc_hd__or3b_1
X_7381_ _7381_/A _7381_/B vssd1 vssd1 vccd1 vccd1 _7382_/B sky130_fd_sc_hd__nand2_1
X_6332_ _6332_/A vssd1 vssd1 vccd1 vccd1 _8528_/D sky130_fd_sc_hd__clkbuf_1
X_6263_ _6082_/A _6249_/A _6263_/S vssd1 vssd1 vccd1 vccd1 _6264_/D sky130_fd_sc_hd__mux2_1
X_5214_ _8558_/Q _5202_/X _5212_/X _5213_/X vssd1 vssd1 vccd1 vccd1 _8483_/D sky130_fd_sc_hd__o211a_1
XFILLER_88_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8002_ _8306_/A _8025_/A vssd1 vssd1 vccd1 vccd1 _8003_/C sky130_fd_sc_hd__nor2_1
X_6194_ _6194_/A _6194_/B vssd1 vssd1 vccd1 vccd1 _6214_/A sky130_fd_sc_hd__xnor2_1
XFILLER_96_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5145_ _4749_/A _5144_/X _4993_/A vssd1 vssd1 vccd1 vccd1 _5160_/D sky130_fd_sc_hd__a21o_1
XFILLER_69_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5076_ _5173_/A _5080_/C _5075_/X vssd1 vssd1 vccd1 vccd1 _5076_/X sky130_fd_sc_hd__or3b_1
XFILLER_56_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8766_ _8766_/A _4356_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[13] sky130_fd_sc_hd__ebufn_8
X_5978_ _5978_/A _5978_/B vssd1 vssd1 vccd1 vccd1 _6106_/A sky130_fd_sc_hd__or2_1
XFILLER_25_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4929_ _4929_/A _4975_/B vssd1 vssd1 vccd1 vccd1 _5159_/B sky130_fd_sc_hd__or2_1
X_8697_ _8697_/A _4276_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[14] sky130_fd_sc_hd__ebufn_8
X_7717_ _7634_/B _7717_/B vssd1 vssd1 vccd1 vccd1 _7758_/A sky130_fd_sc_hd__and2b_1
XFILLER_60_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7648_ _8367_/A _7822_/B vssd1 vssd1 vccd1 vccd1 _7769_/A sky130_fd_sc_hd__nand2_2
XFILLER_20_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7579_ _7607_/A _7583_/A vssd1 vssd1 vccd1 vccd1 _7725_/B sky130_fd_sc_hd__or2_1
XFILLER_85_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8636__52 vssd1 vssd1 vccd1 vccd1 _8636__52/HI _8745_/A sky130_fd_sc_hd__conb_1
XFILLER_78_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6950_ _6991_/A _6932_/B _6949_/Y vssd1 vssd1 vccd1 vccd1 _6952_/A sky130_fd_sc_hd__o21a_1
XFILLER_53_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5901_ _5901_/A vssd1 vssd1 vccd1 vccd1 _6126_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_19_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6881_ _6879_/A _6879_/C _6879_/B vssd1 vssd1 vccd1 vccd1 _6883_/C sky130_fd_sc_hd__a21o_1
X_5832_ _6019_/A _5843_/A _6154_/A vssd1 vssd1 vccd1 vccd1 _5833_/B sky130_fd_sc_hd__o21ba_1
X_8551_ input3/X _8551_/D vssd1 vssd1 vccd1 vccd1 _8551_/Q sky130_fd_sc_hd__dfxtp_1
X_5763_ _5499_/A _5496_/B _5499_/C _5494_/X _5488_/A vssd1 vssd1 vccd1 vccd1 _5943_/A
+ sky130_fd_sc_hd__a311o_2
X_4714_ _7498_/B _4740_/C vssd1 vssd1 vccd1 vccd1 _4738_/B sky130_fd_sc_hd__and2_1
X_7502_ _7500_/X _7505_/A vssd1 vssd1 vccd1 vccd1 _7641_/B sky130_fd_sc_hd__and2b_2
X_8482_ input3/X _8482_/D vssd1 vssd1 vccd1 vccd1 _8482_/Q sky130_fd_sc_hd__dfxtp_1
X_5694_ _5694_/A vssd1 vssd1 vccd1 vccd1 _5805_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4645_ _4649_/B _4645_/B _4645_/C vssd1 vssd1 vccd1 vccd1 _4646_/A sky130_fd_sc_hd__and3b_1
X_7433_ _8575_/Q vssd1 vssd1 vccd1 vccd1 _7539_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7364_ _7365_/A _7365_/B vssd1 vssd1 vccd1 vccd1 _7372_/C sky130_fd_sc_hd__nor2_1
X_4576_ _4576_/A vssd1 vssd1 vccd1 vccd1 _8452_/D sky130_fd_sc_hd__clkbuf_1
X_6315_ _8547_/Q _6315_/B vssd1 vssd1 vccd1 vccd1 _6328_/B sky130_fd_sc_hd__nand2_1
XFILLER_89_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7295_ _7295_/A _7295_/B vssd1 vssd1 vccd1 vccd1 _7301_/A sky130_fd_sc_hd__xnor2_1
X_6246_ _6264_/A _6264_/B _6264_/C _6253_/B vssd1 vssd1 vccd1 vccd1 _6246_/X sky130_fd_sc_hd__or4_1
X_6177_ _6177_/A _6177_/B vssd1 vssd1 vccd1 vccd1 _6228_/A sky130_fd_sc_hd__xor2_1
X_5128_ _5046_/A _5068_/X _5082_/X _5127_/X vssd1 vssd1 vccd1 vccd1 _5128_/X sky130_fd_sc_hd__o31a_1
XFILLER_84_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5059_ _5059_/A vssd1 vssd1 vccd1 vccd1 _5059_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_84_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8749_ _8749_/A _4389_/Y vssd1 vssd1 vccd1 vccd1 io_out[34] sky130_fd_sc_hd__ebufn_8
XFILLER_71_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4430_ _4748_/D vssd1 vssd1 vccd1 vccd1 _4780_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_8_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4361_ _4363_/A vssd1 vssd1 vccd1 vccd1 _4361_/Y sky130_fd_sc_hd__inv_2
X_6100_ _6008_/A _6008_/B _6011_/A vssd1 vssd1 vccd1 vccd1 _6216_/B sky130_fd_sc_hd__o21ai_1
X_4292_ _4295_/A vssd1 vssd1 vccd1 vccd1 _4292_/Y sky130_fd_sc_hd__inv_2
X_7080_ _7085_/A _7085_/B vssd1 vssd1 vccd1 vccd1 _7081_/B sky130_fd_sc_hd__xnor2_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6031_ _6153_/B vssd1 vssd1 vccd1 vccd1 _6033_/A sky130_fd_sc_hd__inv_2
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7982_ _8041_/C _7982_/B vssd1 vssd1 vccd1 vccd1 _7986_/A sky130_fd_sc_hd__xor2_1
XFILLER_26_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6933_ _6996_/A _6996_/B _6996_/C vssd1 vssd1 vccd1 vccd1 _6933_/Y sky130_fd_sc_hd__nand3_2
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6864_ _6863_/A _6863_/C _6863_/B vssd1 vssd1 vccd1 vccd1 _6874_/C sky130_fd_sc_hd__a21o_1
XFILLER_50_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5815_ _5816_/B _5815_/B vssd1 vssd1 vccd1 vccd1 _6061_/B sky130_fd_sc_hd__xnor2_1
XFILLER_34_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6795_ _6795_/A _6795_/B vssd1 vssd1 vccd1 vccd1 _7315_/A sky130_fd_sc_hd__xor2_1
X_8534_ input3/X _8534_/D vssd1 vssd1 vccd1 vccd1 _8534_/Q sky130_fd_sc_hd__dfxtp_1
X_5746_ _5749_/B _5746_/B vssd1 vssd1 vccd1 vccd1 _6057_/A sky130_fd_sc_hd__xnor2_2
XFILLER_41_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8465_ input3/X _8465_/D vssd1 vssd1 vccd1 vccd1 _8465_/Q sky130_fd_sc_hd__dfxtp_1
X_5677_ _5677_/A _5677_/B _5676_/Y vssd1 vssd1 vccd1 vccd1 _6090_/B sky130_fd_sc_hd__or3b_1
X_4628_ _5067_/A vssd1 vssd1 vccd1 vccd1 _5175_/S sky130_fd_sc_hd__clkbuf_2
X_7416_ _8587_/Q vssd1 vssd1 vccd1 vccd1 _7416_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_8396_ _8396_/A vssd1 vssd1 vccd1 vccd1 _8582_/D sky130_fd_sc_hd__clkbuf_1
X_7347_ _7347_/A _7347_/B vssd1 vssd1 vccd1 vccd1 _7347_/Y sky130_fd_sc_hd__xnor2_1
X_4559_ _4561_/B _4568_/B _4559_/C vssd1 vssd1 vccd1 vccd1 _4560_/A sky130_fd_sc_hd__and3b_1
X_7278_ _6891_/A _7276_/X _7277_/X vssd1 vssd1 vccd1 vccd1 _7279_/B sky130_fd_sc_hd__o21ai_1
X_6229_ _6229_/A _6229_/B vssd1 vssd1 vccd1 vccd1 _6230_/B sky130_fd_sc_hd__xnor2_4
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8606__22 vssd1 vssd1 vccd1 vccd1 _8606__22/HI _8701_/A sky130_fd_sc_hd__conb_1
XFILLER_48_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6580_ _6819_/A _6580_/B vssd1 vssd1 vccd1 vccd1 _6581_/B sky130_fd_sc_hd__xor2_2
X_5600_ _6084_/A _5600_/B vssd1 vssd1 vccd1 vccd1 _5673_/A sky130_fd_sc_hd__nand2_1
XFILLER_31_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5531_ _6244_/A _5650_/A vssd1 vssd1 vccd1 vccd1 _5649_/A sky130_fd_sc_hd__nand2_2
X_8250_ _7983_/B _8306_/B _8227_/Y vssd1 vssd1 vccd1 vccd1 _8252_/B sky130_fd_sc_hd__o21a_1
X_7201_ _7201_/A _7201_/B vssd1 vssd1 vccd1 vccd1 _7259_/A sky130_fd_sc_hd__xor2_1
X_5462_ _5459_/A _5459_/B _5437_/A vssd1 vssd1 vccd1 vccd1 _5463_/B sky130_fd_sc_hd__a21oi_1
X_4413_ _7518_/B vssd1 vssd1 vccd1 vccd1 _4698_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5393_ _5417_/A _5404_/B vssd1 vssd1 vccd1 vccd1 _5648_/A sky130_fd_sc_hd__xnor2_4
X_8181_ _8181_/A _8182_/B vssd1 vssd1 vccd1 vccd1 _8194_/B sky130_fd_sc_hd__xnor2_1
X_7132_ _7139_/A _7132_/B vssd1 vssd1 vccd1 vccd1 _7133_/B sky130_fd_sc_hd__xnor2_1
X_4344_ _4345_/A vssd1 vssd1 vccd1 vccd1 _4344_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7063_ _7064_/A _7064_/B _7064_/C vssd1 vssd1 vccd1 vccd1 _7065_/A sky130_fd_sc_hd__a21oi_1
XFILLER_59_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4275_ _4277_/A vssd1 vssd1 vccd1 vccd1 _4275_/Y sky130_fd_sc_hd__inv_2
X_6014_ _6015_/A _6015_/B vssd1 vssd1 vccd1 vccd1 _6014_/X sky130_fd_sc_hd__or2_1
XFILLER_67_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8591__7 vssd1 vssd1 vccd1 vccd1 _8591__7/HI _8686_/A sky130_fd_sc_hd__conb_1
XFILLER_82_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7965_ _8050_/A _7965_/B vssd1 vssd1 vccd1 vccd1 _7966_/B sky130_fd_sc_hd__xnor2_2
XFILLER_82_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6916_ _6916_/A _6916_/B _6916_/C vssd1 vssd1 vccd1 vccd1 _6918_/A sky130_fd_sc_hd__and3_1
X_7896_ _8052_/A _8326_/B vssd1 vssd1 vccd1 vccd1 _7896_/Y sky130_fd_sc_hd__nor2_1
X_6847_ _6854_/A _6847_/B vssd1 vssd1 vccd1 vccd1 _6848_/C sky130_fd_sc_hd__and2_1
XFILLER_50_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6778_ _7026_/A _6778_/B vssd1 vssd1 vccd1 vccd1 _6778_/Y sky130_fd_sc_hd__nand2_1
XFILLER_10_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8517_ input3/X _8517_/D vssd1 vssd1 vccd1 vccd1 _8517_/Q sky130_fd_sc_hd__dfxtp_1
X_5729_ _6188_/B _6025_/A vssd1 vssd1 vccd1 vccd1 _5734_/A sky130_fd_sc_hd__or2_1
X_8448_ input3/X _8448_/D vssd1 vssd1 vccd1 vccd1 _8448_/Q sky130_fd_sc_hd__dfxtp_1
X_8379_ _8373_/X _8378_/X _6261_/X _8578_/Q vssd1 vssd1 vccd1 vccd1 _8578_/D sky130_fd_sc_hd__o2bb2a_1
XFILLER_2_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4962_ _5074_/A _5116_/B vssd1 vssd1 vccd1 vccd1 _4962_/X sky130_fd_sc_hd__or2_1
X_7750_ _7750_/A _7750_/B _7750_/C vssd1 vssd1 vccd1 vccd1 _7751_/B sky130_fd_sc_hd__nand3_1
X_4893_ _4893_/A _5156_/A _4862_/A vssd1 vssd1 vccd1 vccd1 _4893_/X sky130_fd_sc_hd__or3b_1
X_6701_ _6698_/A _6698_/B _6698_/C _6725_/A vssd1 vssd1 vccd1 vccd1 _6727_/A sky130_fd_sc_hd__a31o_1
X_7681_ _8099_/A _7681_/B vssd1 vssd1 vccd1 vccd1 _8101_/C sky130_fd_sc_hd__nand2_1
XFILLER_32_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6632_ _6632_/A _7043_/B _6810_/A vssd1 vssd1 vccd1 vccd1 _6755_/A sky130_fd_sc_hd__or3_1
XFILLER_32_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6563_ _6563_/A _6563_/B vssd1 vssd1 vccd1 vccd1 _6652_/B sky130_fd_sc_hd__nor2_1
X_6494_ _8467_/Q _8550_/Q vssd1 vssd1 vccd1 vccd1 _6501_/A sky130_fd_sc_hd__or2b_1
X_8302_ _8302_/A _8302_/B vssd1 vssd1 vccd1 vccd1 _8302_/Y sky130_fd_sc_hd__nand2_1
X_5514_ _5940_/A _6026_/A vssd1 vssd1 vccd1 vccd1 _5515_/C sky130_fd_sc_hd__nand2_1
X_8233_ _8233_/A _8233_/B _8233_/C vssd1 vssd1 vccd1 vccd1 _8234_/B sky130_fd_sc_hd__nor3_1
X_5445_ _5445_/A _5445_/B vssd1 vssd1 vccd1 vccd1 _5609_/A sky130_fd_sc_hd__xor2_1
X_8164_ _8165_/A _8165_/B _8165_/C vssd1 vssd1 vccd1 vccd1 _8166_/A sky130_fd_sc_hd__o21a_1
X_7115_ _7134_/A _7134_/B vssd1 vssd1 vccd1 vccd1 _7161_/A sky130_fd_sc_hd__xor2_1
X_5376_ _5651_/A vssd1 vssd1 vccd1 vccd1 _5705_/A sky130_fd_sc_hd__clkbuf_2
X_4327_ _4327_/A vssd1 vssd1 vccd1 vccd1 _4332_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_86_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8095_ _7697_/A _8366_/A _8105_/B vssd1 vssd1 vccd1 vccd1 _8104_/A sky130_fd_sc_hd__a21o_1
X_4258_ _4382_/A vssd1 vssd1 vccd1 vccd1 _4390_/A sky130_fd_sc_hd__buf_6
X_7046_ _7101_/A _7102_/A _7036_/X _7040_/Y _7033_/X vssd1 vssd1 vccd1 vccd1 _7099_/A
+ sky130_fd_sc_hd__o2111ai_2
XFILLER_74_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8597__13 vssd1 vssd1 vccd1 vccd1 _8597__13/HI _8692_/A sky130_fd_sc_hd__conb_1
XFILLER_82_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7948_ _7621_/B _8063_/B _7947_/X vssd1 vssd1 vccd1 vccd1 _7949_/B sky130_fd_sc_hd__o21ba_1
XFILLER_42_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7879_ _7877_/X _7867_/B _7878_/X vssd1 vssd1 vccd1 vccd1 _7904_/A sky130_fd_sc_hd__o21bai_4
XFILLER_10_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5230_ _8486_/Q _5230_/B vssd1 vssd1 vccd1 vccd1 _5231_/A sky130_fd_sc_hd__and2b_1
XFILLER_5_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5161_ _4886_/A _5071_/A _5012_/A vssd1 vssd1 vccd1 vccd1 _5164_/C sky130_fd_sc_hd__o21a_1
XFILLER_69_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5092_ _5092_/A _5092_/B _5092_/C _5092_/D vssd1 vssd1 vccd1 vccd1 _5092_/X sky130_fd_sc_hd__or4_1
XFILLER_96_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8681__97 vssd1 vssd1 vccd1 vccd1 _8681__97/HI _8790_/A sky130_fd_sc_hd__conb_1
XFILLER_52_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8782_ _8782_/A _4377_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[29] sky130_fd_sc_hd__ebufn_8
XFILLER_64_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5994_ _5994_/A _5994_/B vssd1 vssd1 vccd1 vccd1 _6046_/A sky130_fd_sc_hd__xnor2_1
X_7802_ _7802_/A _7802_/B vssd1 vssd1 vccd1 vccd1 _7932_/A sky130_fd_sc_hd__and2_1
X_4945_ _4945_/A _4945_/B vssd1 vssd1 vccd1 vccd1 _4945_/Y sky130_fd_sc_hd__nand2_1
X_7733_ _7733_/A _7888_/B vssd1 vssd1 vccd1 vccd1 _7746_/A sky130_fd_sc_hd__or2_1
X_4876_ _8455_/Q _5026_/A vssd1 vssd1 vccd1 vccd1 _5156_/B sky130_fd_sc_hd__or2_1
X_7664_ _7664_/A _7664_/B vssd1 vssd1 vccd1 vccd1 _7665_/B sky130_fd_sc_hd__or2_1
X_6615_ _6640_/A _6622_/B _7032_/B _6736_/B vssd1 vssd1 vccd1 vccd1 _6616_/C sky130_fd_sc_hd__or4_1
X_7595_ _7725_/A vssd1 vssd1 vccd1 vccd1 _7731_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6546_ _6603_/A _8470_/Q _6500_/A _6500_/B _6499_/A vssd1 vssd1 vccd1 vccd1 _6596_/B
+ sky130_fd_sc_hd__a221o_1
X_6477_ _8563_/Q _8459_/Q vssd1 vssd1 vccd1 vccd1 _6479_/A sky130_fd_sc_hd__and2b_1
X_5428_ _5429_/A _5429_/B _5427_/Y _5537_/B vssd1 vssd1 vccd1 vccd1 _5557_/A sky130_fd_sc_hd__a22oi_2
X_8216_ _8202_/A _8204_/A _8192_/B vssd1 vssd1 vccd1 vccd1 _8216_/X sky130_fd_sc_hd__o21a_1
X_8147_ _8147_/A _8147_/B vssd1 vssd1 vccd1 vccd1 _8154_/A sky130_fd_sc_hd__nor2_1
X_5359_ _5360_/A _5359_/B vssd1 vssd1 vccd1 vccd1 _5362_/C sky130_fd_sc_hd__nand2_1
XINSDIODE2_2 _7201_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8078_ _8078_/A _8078_/B vssd1 vssd1 vccd1 vccd1 _8088_/B sky130_fd_sc_hd__xnor2_2
X_7029_ _7272_/B _7272_/C vssd1 vssd1 vccd1 vccd1 _7030_/B sky130_fd_sc_hd__nand2_1
XFILLER_47_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4730_ _5040_/B _5153_/B vssd1 vssd1 vccd1 vccd1 _5169_/A sky130_fd_sc_hd__or2_2
XFILLER_14_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4661_ _7478_/A _4661_/B vssd1 vssd1 vccd1 vccd1 _4661_/X sky130_fd_sc_hd__or2_1
XFILLER_9_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7380_ _7380_/A _8548_/Q vssd1 vssd1 vccd1 vccd1 _7381_/B sky130_fd_sc_hd__or2b_1
X_6400_ _8548_/Q vssd1 vssd1 vccd1 vccd1 _7390_/A sky130_fd_sc_hd__clkbuf_1
X_4592_ _4592_/A _4663_/A vssd1 vssd1 vccd1 vccd1 _4619_/B sky130_fd_sc_hd__nand2_1
X_6331_ _6322_/A _6331_/B _6331_/C vssd1 vssd1 vccd1 vccd1 _6332_/A sky130_fd_sc_hd__and3b_1
X_6262_ _6251_/X _6260_/X _6261_/X _8518_/Q vssd1 vssd1 vccd1 vccd1 _8518_/D sky130_fd_sc_hd__o2bb2a_1
XFILLER_88_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6193_ _6193_/A _6193_/B vssd1 vssd1 vccd1 vccd1 _6194_/B sky130_fd_sc_hd__xnor2_1
X_8001_ _8105_/A vssd1 vssd1 vccd1 vccd1 _8306_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5213_ _8419_/A vssd1 vssd1 vccd1 vccd1 _5213_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_69_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5144_ _4737_/A _5144_/B _5144_/C vssd1 vssd1 vccd1 vccd1 _5144_/X sky130_fd_sc_hd__and3b_1
XFILLER_57_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5075_ _5160_/A _5073_/Y _5074_/Y _4963_/X _5080_/A vssd1 vssd1 vccd1 vccd1 _5075_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_84_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8765_ _8765_/A _4354_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[12] sky130_fd_sc_hd__ebufn_8
XFILLER_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5977_ _5861_/C _5975_/X _5976_/X vssd1 vssd1 vccd1 vccd1 _6104_/A sky130_fd_sc_hd__o21ai_2
XFILLER_40_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4928_ _5012_/A _5160_/C _5064_/C _4927_/X vssd1 vssd1 vccd1 vccd1 _4930_/B sky130_fd_sc_hd__o31a_1
X_8696_ _8696_/A _4275_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[13] sky130_fd_sc_hd__ebufn_8
XFILLER_33_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7716_ _8207_/A _7716_/B vssd1 vssd1 vccd1 vccd1 _7792_/A sky130_fd_sc_hd__nand2_1
XFILLER_40_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7647_ _7647_/A _7647_/B vssd1 vssd1 vccd1 vccd1 _7822_/B sky130_fd_sc_hd__xnor2_4
X_4859_ _5036_/A _5058_/B _5138_/C vssd1 vssd1 vccd1 vccd1 _4859_/X sky130_fd_sc_hd__or3_1
X_7578_ _7606_/A _7606_/B vssd1 vssd1 vccd1 vccd1 _7583_/A sky130_fd_sc_hd__xnor2_2
X_6529_ _6507_/A _6557_/A _6531_/A vssd1 vssd1 vccd1 vccd1 _6761_/A sky130_fd_sc_hd__mux2_2
XFILLER_4_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8651__67 vssd1 vssd1 vccd1 vccd1 _8651__67/HI _8760_/A sky130_fd_sc_hd__conb_1
XFILLER_38_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5900_ _5900_/A _5900_/B vssd1 vssd1 vccd1 vccd1 _6210_/A sky130_fd_sc_hd__nand2_1
XFILLER_19_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6880_ _6880_/A _6880_/B _6880_/C vssd1 vssd1 vccd1 vccd1 _6883_/B sky130_fd_sc_hd__nand3_1
XFILLER_34_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5831_ _5831_/A _6025_/B vssd1 vssd1 vccd1 vccd1 _6154_/A sky130_fd_sc_hd__nor2_2
XFILLER_34_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8550_ input3/X _8550_/D vssd1 vssd1 vccd1 vccd1 _8550_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_61_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5762_ _6188_/B _5825_/B _5825_/C _5838_/A _5738_/A vssd1 vssd1 vccd1 vccd1 _5765_/B
+ sky130_fd_sc_hd__o32ai_4
X_4713_ _4713_/A _4740_/C vssd1 vssd1 vccd1 vccd1 _4737_/A sky130_fd_sc_hd__nor2_1
X_7501_ _7501_/A _7501_/B vssd1 vssd1 vccd1 vccd1 _7505_/A sky130_fd_sc_hd__nand2_1
X_8481_ input3/X _8481_/D vssd1 vssd1 vccd1 vccd1 _8481_/Q sky130_fd_sc_hd__dfxtp_1
X_5693_ _5811_/A _5811_/B vssd1 vssd1 vccd1 vccd1 _5698_/A sky130_fd_sc_hd__xnor2_1
XFILLER_30_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4644_ _4620_/A _4639_/A _5178_/B vssd1 vssd1 vccd1 vccd1 _4645_/C sky130_fd_sc_hd__a21o_1
X_7432_ _7482_/B vssd1 vssd1 vccd1 vccd1 _7481_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_7363_ _6472_/X _8557_/Q _7357_/X _7362_/X vssd1 vssd1 vccd1 vccd1 _8557_/D sky130_fd_sc_hd__o22a_1
X_4575_ _4575_/A _4575_/B _4575_/C vssd1 vssd1 vccd1 vccd1 _4576_/A sky130_fd_sc_hd__and3_1
XFILLER_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6314_ _8545_/Q _6313_/X _8546_/Q vssd1 vssd1 vccd1 vccd1 _6315_/B sky130_fd_sc_hd__a21o_1
X_7294_ _7323_/A _7294_/B vssd1 vssd1 vccd1 vccd1 _7295_/B sky130_fd_sc_hd__nor2_1
X_6245_ _6247_/A _6243_/Y _6244_/X _5455_/B vssd1 vssd1 vccd1 vccd1 _6253_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_39_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6176_ _5860_/A _6126_/A _6184_/B _5918_/C vssd1 vssd1 vccd1 vccd1 _6177_/B sky130_fd_sc_hd__o22a_1
X_5127_ _4863_/X _5098_/X _5109_/X _5126_/X _5046_/Y vssd1 vssd1 vccd1 vccd1 _5127_/X
+ sky130_fd_sc_hd__a311o_1
X_5058_ _5099_/B _5058_/B _5058_/C vssd1 vssd1 vccd1 vccd1 _5058_/X sky130_fd_sc_hd__or3_1
XFILLER_84_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8748_ _8748_/A _4338_/Y vssd1 vssd1 vccd1 vccd1 io_out[33] sky130_fd_sc_hd__ebufn_8
XFILLER_52_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4360_ _4363_/A vssd1 vssd1 vccd1 vccd1 _4360_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4291_ _4295_/A vssd1 vssd1 vccd1 vccd1 _4291_/Y sky130_fd_sc_hd__inv_2
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6030_ _6030_/A _6030_/B vssd1 vssd1 vccd1 vccd1 _6036_/A sky130_fd_sc_hd__xor2_2
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7981_ _7813_/A _7925_/B _8120_/A _7980_/Y vssd1 vssd1 vccd1 vccd1 _7982_/B sky130_fd_sc_hd__a31o_1
X_6932_ _6991_/A _6932_/B vssd1 vssd1 vccd1 vccd1 _6996_/C sky130_fd_sc_hd__xor2_2
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6863_ _6863_/A _6863_/B _6863_/C vssd1 vssd1 vccd1 vccd1 _6874_/B sky130_fd_sc_hd__nand3_1
X_5814_ _5814_/A _5814_/B vssd1 vssd1 vccd1 vccd1 _5815_/B sky130_fd_sc_hd__xnor2_1
XFILLER_22_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6794_ _6794_/A _6794_/B vssd1 vssd1 vccd1 vccd1 _6795_/B sky130_fd_sc_hd__nor2_1
XFILLER_22_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8533_ input3/X _8533_/D vssd1 vssd1 vccd1 vccd1 _8533_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5745_ _5745_/A _5745_/B vssd1 vssd1 vccd1 vccd1 _5746_/B sky130_fd_sc_hd__xnor2_1
X_8464_ input3/X _8464_/D vssd1 vssd1 vccd1 vccd1 _8464_/Q sky130_fd_sc_hd__dfxtp_1
X_5676_ _6070_/B _5676_/B vssd1 vssd1 vccd1 vccd1 _5676_/Y sky130_fd_sc_hd__nand2_1
X_4627_ _4862_/A _4862_/B vssd1 vssd1 vccd1 vccd1 _5067_/A sky130_fd_sc_hd__or2_1
X_7415_ _8585_/Q vssd1 vssd1 vccd1 vccd1 _8428_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_8395_ _8403_/A _8395_/B vssd1 vssd1 vccd1 vccd1 _8396_/A sky130_fd_sc_hd__and2_1
X_7346_ _7338_/A _7341_/B _7338_/C _7345_/Y vssd1 vssd1 vccd1 vccd1 _7347_/B sky130_fd_sc_hd__a31o_1
X_4558_ _8446_/Q _8445_/Q _4552_/B _8447_/Q vssd1 vssd1 vccd1 vccd1 _4559_/C sky130_fd_sc_hd__a31o_1
X_4489_ _8478_/Q _4491_/B vssd1 vssd1 vccd1 vccd1 _4490_/A sky130_fd_sc_hd__and2_1
XFILLER_89_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7277_ _7277_/A _6890_/A vssd1 vssd1 vccd1 vccd1 _7277_/X sky130_fd_sc_hd__or2b_1
XFILLER_89_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6228_ _6228_/A _6228_/B vssd1 vssd1 vccd1 vccd1 _6229_/B sky130_fd_sc_hd__xnor2_2
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6159_ _6160_/A _6160_/B vssd1 vssd1 vccd1 vccd1 _6159_/X sky130_fd_sc_hd__and2_1
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8621__37 vssd1 vssd1 vccd1 vccd1 _8621__37/HI _8716_/A sky130_fd_sc_hd__conb_1
XFILLER_91_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5530_ _5530_/A _5530_/B vssd1 vssd1 vccd1 vccd1 _5650_/A sky130_fd_sc_hd__xnor2_2
XFILLER_8_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5461_ _5461_/A _5461_/B vssd1 vssd1 vccd1 vccd1 _5463_/A sky130_fd_sc_hd__nand2_1
X_7200_ _7200_/A _7200_/B _7200_/C vssd1 vssd1 vccd1 vccd1 _7341_/B sky130_fd_sc_hd__nand3_2
X_4412_ _8471_/Q vssd1 vssd1 vccd1 vccd1 _7518_/B sky130_fd_sc_hd__buf_2
XFILLER_8_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5392_ _5686_/A vssd1 vssd1 vccd1 vccd1 _5685_/A sky130_fd_sc_hd__clkbuf_2
X_8180_ _8180_/A _8180_/B vssd1 vssd1 vccd1 vccd1 _8182_/B sky130_fd_sc_hd__xor2_1
X_7131_ _7131_/A _7131_/B vssd1 vssd1 vccd1 vccd1 _7132_/B sky130_fd_sc_hd__xor2_1
X_4343_ _4345_/A vssd1 vssd1 vccd1 vccd1 _4343_/Y sky130_fd_sc_hd__inv_2
X_7062_ _7062_/A _7062_/B vssd1 vssd1 vccd1 vccd1 _7064_/C sky130_fd_sc_hd__xnor2_1
X_4274_ _4277_/A vssd1 vssd1 vccd1 vccd1 _4274_/Y sky130_fd_sc_hd__inv_2
X_6013_ _5955_/A _6013_/B vssd1 vssd1 vccd1 vccd1 _6042_/B sky130_fd_sc_hd__and2b_1
XFILLER_39_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7964_ _7964_/A _7964_/B vssd1 vssd1 vccd1 vccd1 _7965_/B sky130_fd_sc_hd__xor2_1
XFILLER_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6915_ _6745_/B _6643_/C _6739_/A _6586_/A vssd1 vssd1 vccd1 vccd1 _6916_/C sky130_fd_sc_hd__a31o_1
X_7895_ _8147_/B vssd1 vssd1 vccd1 vccd1 _8326_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_35_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6846_ _6893_/A _6846_/B vssd1 vssd1 vccd1 vccd1 _6847_/B sky130_fd_sc_hd__or2_1
XFILLER_22_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6777_ _6777_/A _6777_/B vssd1 vssd1 vccd1 vccd1 _6791_/B sky130_fd_sc_hd__and2_1
X_8516_ input3/X _8516_/D vssd1 vssd1 vccd1 vccd1 _8516_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5728_ _5758_/A _5758_/B vssd1 vssd1 vccd1 vccd1 _5735_/A sky130_fd_sc_hd__xnor2_1
X_8447_ input3/X _8447_/D vssd1 vssd1 vccd1 vccd1 _8447_/Q sky130_fd_sc_hd__dfxtp_1
X_5659_ _5659_/A _5659_/B vssd1 vssd1 vccd1 vccd1 _5660_/B sky130_fd_sc_hd__and2_1
X_8378_ _8385_/A _8385_/B _8385_/C _8378_/D vssd1 vssd1 vccd1 vccd1 _8378_/X sky130_fd_sc_hd__or4_1
X_7329_ _7329_/A _7329_/B vssd1 vssd1 vccd1 vccd1 _7330_/B sky130_fd_sc_hd__xnor2_1
XFILLER_93_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4961_ _5117_/A _5025_/A vssd1 vssd1 vccd1 vccd1 _5116_/B sky130_fd_sc_hd__or2_2
XFILLER_17_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4892_ _4987_/A _4874_/X _5156_/B _4891_/X vssd1 vssd1 vccd1 vccd1 _4893_/A sky130_fd_sc_hd__o31a_1
X_6700_ _6700_/A _6700_/B _6700_/C vssd1 vssd1 vccd1 vccd1 _6725_/A sky130_fd_sc_hd__and3_1
XFILLER_32_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7680_ _7680_/A _7680_/B vssd1 vssd1 vccd1 vccd1 _7681_/B sky130_fd_sc_hd__xor2_1
X_6631_ _6736_/A vssd1 vssd1 vccd1 vccd1 _6810_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_32_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6562_ _7575_/B _6562_/B vssd1 vssd1 vccd1 vccd1 _6563_/A sky130_fd_sc_hd__and2b_1
X_8301_ _8240_/A _8240_/B _8241_/B _8241_/A vssd1 vssd1 vccd1 vccd1 _8311_/A sky130_fd_sc_hd__a2bb2o_1
X_6493_ _6501_/B _7233_/A vssd1 vssd1 vccd1 vccd1 _6508_/C sky130_fd_sc_hd__or2b_1
X_5513_ _5764_/B _5764_/C vssd1 vssd1 vccd1 vccd1 _6026_/A sky130_fd_sc_hd__or2_2
X_8232_ _8233_/A _8233_/B _8233_/C vssd1 vssd1 vccd1 vccd1 _8234_/A sky130_fd_sc_hd__o21a_1
X_5444_ _5461_/A _5444_/B vssd1 vssd1 vccd1 vccd1 _5445_/B sky130_fd_sc_hd__nand2_1
X_8163_ _8163_/A _8163_/B vssd1 vssd1 vccd1 vccd1 _8165_/C sky130_fd_sc_hd__xor2_1
X_7114_ _7114_/A _7114_/B vssd1 vssd1 vccd1 vccd1 _7134_/B sky130_fd_sc_hd__xnor2_1
X_5375_ _5417_/A _5417_/B vssd1 vssd1 vccd1 vccd1 _5651_/A sky130_fd_sc_hd__and2_1
X_4326_ _4326_/A vssd1 vssd1 vccd1 vccd1 _4326_/Y sky130_fd_sc_hd__inv_2
X_8094_ _8023_/A _8023_/B _8028_/B _8093_/Y vssd1 vssd1 vccd1 vccd1 _8238_/B sky130_fd_sc_hd__a31o_1
X_4257_ input1/X vssd1 vssd1 vccd1 vccd1 _4382_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_86_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7045_ _7105_/A _7045_/B vssd1 vssd1 vccd1 vccd1 _7099_/C sky130_fd_sc_hd__xor2_1
XFILLER_74_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7947_ _7731_/A _7885_/B _7885_/C _7950_/A _7620_/A vssd1 vssd1 vccd1 vccd1 _7947_/X
+ sky130_fd_sc_hd__o32a_1
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7878_ _7877_/B _7878_/B vssd1 vssd1 vccd1 vccd1 _7878_/X sky130_fd_sc_hd__and2b_1
X_6829_ _6829_/A vssd1 vssd1 vccd1 vccd1 _6874_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_10_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5160_ _5160_/A _5173_/A _5160_/C _5160_/D vssd1 vssd1 vccd1 vccd1 _5160_/X sky130_fd_sc_hd__or4_1
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5091_ _5091_/A _5118_/B vssd1 vssd1 vccd1 vccd1 _5091_/X sky130_fd_sc_hd__or2_1
XFILLER_68_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8781_ _8781_/A _4375_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[28] sky130_fd_sc_hd__ebufn_8
XFILLER_52_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7801_ _8372_/A _8381_/A _8372_/B vssd1 vssd1 vccd1 vccd1 _8385_/A sky130_fd_sc_hd__a21oi_1
X_5993_ _5993_/A _5993_/B vssd1 vssd1 vccd1 vccd1 _5994_/B sky130_fd_sc_hd__xor2_2
XFILLER_91_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4944_ _4944_/A _4944_/B vssd1 vssd1 vccd1 vccd1 _4945_/B sky130_fd_sc_hd__or2_1
XFILLER_52_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7732_ _7618_/A _7615_/B _7618_/C _7613_/X vssd1 vssd1 vccd1 vccd1 _7888_/B sky130_fd_sc_hd__a31o_1
X_4875_ _4899_/A _4875_/B vssd1 vssd1 vccd1 vccd1 _5026_/A sky130_fd_sc_hd__nor2_1
X_7663_ _7664_/A _7664_/B vssd1 vssd1 vccd1 vccd1 _7665_/A sky130_fd_sc_hd__nand2_1
X_6614_ _6614_/A vssd1 vssd1 vccd1 vccd1 _7032_/B sky130_fd_sc_hd__clkbuf_2
X_7594_ _7594_/A _7594_/B vssd1 vssd1 vccd1 vccd1 _7725_/A sky130_fd_sc_hd__nand2_1
X_6545_ _6603_/A _8470_/Q vssd1 vssd1 vccd1 vccd1 _6604_/A sky130_fd_sc_hd__or2_1
XFILLER_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6476_ _6486_/A _6486_/B _6475_/X vssd1 vssd1 vccd1 vccd1 _6999_/A sky130_fd_sc_hd__a21o_2
X_8215_ _8361_/A _8361_/B _8212_/X _8214_/X vssd1 vssd1 vccd1 vccd1 _8355_/B sky130_fd_sc_hd__a31o_1
X_8657__73 vssd1 vssd1 vccd1 vccd1 _8657__73/HI _8766_/A sky130_fd_sc_hd__conb_1
X_5427_ _5522_/A _5427_/B vssd1 vssd1 vccd1 vccd1 _5427_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_87_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5358_ _5333_/A _5356_/X _5367_/S _5332_/X _5366_/A vssd1 vssd1 vccd1 vccd1 _8513_/D
+ sky130_fd_sc_hd__a32o_1
X_8146_ _8146_/A _8146_/B vssd1 vssd1 vccd1 vccd1 _8148_/A sky130_fd_sc_hd__nor2_2
X_4309_ _4327_/A vssd1 vssd1 vccd1 vccd1 _4314_/A sky130_fd_sc_hd__clkbuf_2
XINSDIODE2_3 _7201_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8077_ _8077_/A _8116_/B vssd1 vssd1 vccd1 vccd1 _8078_/B sky130_fd_sc_hd__xnor2_1
X_7028_ _7146_/A _7272_/B _7028_/C vssd1 vssd1 vccd1 vccd1 _7272_/C sky130_fd_sc_hd__nand3_1
XFILLER_87_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5289_ _8504_/Q _5290_/B vssd1 vssd1 vccd1 vccd1 _5291_/B sky130_fd_sc_hd__or2_1
XFILLER_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4660_ _4754_/B _4663_/B vssd1 vssd1 vccd1 vccd1 _4661_/B sky130_fd_sc_hd__nor2_1
XFILLER_80_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4591_ _7766_/B _4706_/A _4591_/C _4747_/A vssd1 vssd1 vccd1 vccd1 _4663_/A sky130_fd_sc_hd__or4_2
X_6330_ _8528_/Q _8527_/Q vssd1 vssd1 vccd1 vccd1 _6331_/C sky130_fd_sc_hd__nand2_1
X_6261_ _7412_/A vssd1 vssd1 vccd1 vccd1 _6261_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5212_ _8483_/Q _5217_/B vssd1 vssd1 vccd1 vccd1 _5212_/X sky130_fd_sc_hd__or2_1
X_6192_ _6192_/A _6192_/B vssd1 vssd1 vccd1 vccd1 _6193_/B sky130_fd_sc_hd__xnor2_1
X_8000_ _8241_/A _8022_/B vssd1 vssd1 vccd1 vccd1 _8003_/B sky130_fd_sc_hd__xor2_1
XFILLER_96_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5143_ _5099_/B _5030_/B _5142_/X _5153_/B _4839_/A vssd1 vssd1 vccd1 vccd1 _5146_/C
+ sky130_fd_sc_hd__o32a_1
X_5074_ _5074_/A _5074_/B vssd1 vssd1 vccd1 vccd1 _5074_/Y sky130_fd_sc_hd__nor2_1
XFILLER_84_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8764_ _8764_/A _4351_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[11] sky130_fd_sc_hd__ebufn_8
XFILLER_52_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5976_ _5976_/A _6126_/B vssd1 vssd1 vccd1 vccd1 _5976_/X sky130_fd_sc_hd__or2_1
X_4927_ _5019_/A _5171_/B _4985_/A _5012_/C vssd1 vssd1 vccd1 vccd1 _4927_/X sky130_fd_sc_hd__or4_1
X_8695_ _8695_/A _4274_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[12] sky130_fd_sc_hd__ebufn_8
X_7715_ _7715_/A _7715_/B vssd1 vssd1 vccd1 vccd1 _7716_/B sky130_fd_sc_hd__nand2_1
X_4858_ _5099_/C vssd1 vssd1 vccd1 vccd1 _5058_/B sky130_fd_sc_hd__clkbuf_2
X_7646_ _7542_/A _7539_/Y _7542_/B _7540_/A vssd1 vssd1 vccd1 vccd1 _7647_/B sky130_fd_sc_hd__a31o_2
X_4789_ _4818_/B vssd1 vssd1 vccd1 vccd1 _4953_/B sky130_fd_sc_hd__buf_2
X_7577_ _7574_/A _7574_/B _7556_/A vssd1 vssd1 vccd1 vccd1 _7606_/B sky130_fd_sc_hd__a21oi_2
X_6528_ _6513_/X _6649_/B _6524_/A _6512_/A _6481_/A vssd1 vssd1 vccd1 vccd1 _6531_/A
+ sky130_fd_sc_hd__a311o_1
XFILLER_69_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6459_ _6459_/A _6466_/A _6466_/B _6459_/D vssd1 vssd1 vccd1 vccd1 _6459_/Y sky130_fd_sc_hd__nand4_1
XFILLER_0_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8129_ _8129_/A _8129_/B vssd1 vssd1 vccd1 vccd1 _8131_/B sky130_fd_sc_hd__xor2_1
XFILLER_87_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5830_ _5765_/A _5765_/B _5765_/C vssd1 vssd1 vccd1 vccd1 _5843_/A sky130_fd_sc_hd__a21bo_1
XFILLER_22_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5761_ _5767_/B vssd1 vssd1 vccd1 vccd1 _5838_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_91_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8480_ input3/X _8480_/D vssd1 vssd1 vccd1 vccd1 _8480_/Q sky130_fd_sc_hd__dfxtp_1
X_4712_ _8466_/Q _8465_/Q _7494_/B vssd1 vssd1 vccd1 vccd1 _4740_/C sky130_fd_sc_hd__o21a_1
X_7500_ _8572_/Q _8469_/Q vssd1 vssd1 vccd1 vccd1 _7500_/X sky130_fd_sc_hd__and2b_1
X_7431_ _8569_/Q vssd1 vssd1 vccd1 vccd1 _7482_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_5692_ _5809_/A _5692_/B vssd1 vssd1 vccd1 vccd1 _5811_/B sky130_fd_sc_hd__and2_1
XFILLER_30_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4643_ _4643_/A _4711_/B vssd1 vssd1 vccd1 vccd1 _4649_/B sky130_fd_sc_hd__nor2_1
X_7362_ _7356_/A _7356_/B _7356_/C _7361_/X _7478_/A vssd1 vssd1 vccd1 vccd1 _7362_/X
+ sky130_fd_sc_hd__a41o_1
X_4574_ _8452_/Q _4574_/B vssd1 vssd1 vccd1 vccd1 _4575_/C sky130_fd_sc_hd__nand2_1
X_6313_ _8542_/Q _6380_/B _6320_/A _6312_/X _8544_/Q vssd1 vssd1 vccd1 vccd1 _6313_/X
+ sky130_fd_sc_hd__a221o_1
X_7293_ _7293_/A _7293_/B vssd1 vssd1 vccd1 vccd1 _7295_/A sky130_fd_sc_hd__or2_1
X_6244_ _6244_/A _6244_/B _5466_/A vssd1 vssd1 vccd1 vccd1 _6244_/X sky130_fd_sc_hd__or3b_1
X_8627__43 vssd1 vssd1 vccd1 vccd1 _8627__43/HI _8722_/A sky130_fd_sc_hd__conb_1
X_6175_ _6168_/A _6168_/B _6173_/X _6174_/Y vssd1 vssd1 vccd1 vccd1 _6229_/A sky130_fd_sc_hd__a211o_2
X_5126_ _5109_/B _5120_/X _5125_/X _5175_/S vssd1 vssd1 vccd1 vccd1 _5126_/X sky130_fd_sc_hd__o211a_1
X_5057_ _5089_/A _5057_/B vssd1 vssd1 vccd1 vccd1 _5057_/X sky130_fd_sc_hd__or2_1
XFILLER_57_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8747_ _8747_/A _4337_/Y vssd1 vssd1 vccd1 vccd1 io_out[32] sky130_fd_sc_hd__ebufn_8
XFILLER_80_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5959_ _5959_/A _5959_/B vssd1 vssd1 vccd1 vccd1 _5963_/B sky130_fd_sc_hd__xnor2_1
XFILLER_40_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7629_ _8070_/A vssd1 vssd1 vccd1 vccd1 _7756_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4290_ _4296_/A vssd1 vssd1 vccd1 vccd1 _4295_/A sky130_fd_sc_hd__clkbuf_2
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7980_ _7984_/A _7921_/B _7984_/C vssd1 vssd1 vccd1 vccd1 _7980_/Y sky130_fd_sc_hd__a21boi_1
X_6931_ _6949_/A _6949_/B vssd1 vssd1 vccd1 vccd1 _6932_/B sky130_fd_sc_hd__xnor2_2
XFILLER_35_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6862_ _6862_/A _6862_/B vssd1 vssd1 vccd1 vccd1 _7319_/A sky130_fd_sc_hd__xnor2_2
XFILLER_62_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5813_ _5813_/A _5813_/B vssd1 vssd1 vccd1 vccd1 _5814_/B sky130_fd_sc_hd__xor2_1
XFILLER_34_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6793_ _6792_/B _6792_/C _7310_/S vssd1 vssd1 vccd1 vccd1 _6794_/B sky130_fd_sc_hd__a21oi_1
X_8532_ input3/X _8532_/D vssd1 vssd1 vccd1 vccd1 _8532_/Q sky130_fd_sc_hd__dfxtp_1
X_5744_ _5744_/A _5751_/B vssd1 vssd1 vccd1 vccd1 _5745_/B sky130_fd_sc_hd__xnor2_1
X_8463_ input3/X _8463_/D vssd1 vssd1 vccd1 vccd1 _8463_/Q sky130_fd_sc_hd__dfxtp_2
X_5675_ _5677_/A _5677_/B _6070_/B _5676_/B vssd1 vssd1 vccd1 vccd1 _6087_/A sky130_fd_sc_hd__o211a_1
X_4626_ _4626_/A _4626_/B vssd1 vssd1 vccd1 vccd1 _4862_/B sky130_fd_sc_hd__nor2_2
X_7414_ _8586_/Q vssd1 vssd1 vccd1 vccd1 _8423_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_8394_ _8393_/Y _8391_/A _8418_/S vssd1 vssd1 vccd1 vccd1 _8395_/B sky130_fd_sc_hd__mux2_1
X_7345_ _7345_/A _7345_/B _7345_/C vssd1 vssd1 vccd1 vccd1 _7345_/Y sky130_fd_sc_hd__nor3_1
X_4557_ _8446_/Q _8447_/Q _4557_/C vssd1 vssd1 vccd1 vccd1 _4561_/B sky130_fd_sc_hd__and3_1
X_4488_ _4488_/A vssd1 vssd1 vccd1 vccd1 _8739_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7276_ _6890_/A _7277_/A vssd1 vssd1 vccd1 vccd1 _7276_/X sky130_fd_sc_hd__and2b_1
XFILLER_1_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6227_ _6227_/A _6227_/B vssd1 vssd1 vccd1 vccd1 _6228_/B sky130_fd_sc_hd__xnor2_1
XFILLER_85_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6158_ _6158_/A _6158_/B vssd1 vssd1 vccd1 vccd1 _6162_/A sky130_fd_sc_hd__xor2_1
X_5109_ _5109_/A _5109_/B _5109_/C _5109_/D vssd1 vssd1 vccd1 vccd1 _5109_/X sky130_fd_sc_hd__or4_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6089_ _6233_/A _6233_/B vssd1 vssd1 vccd1 vccd1 _6089_/X sky130_fd_sc_hd__or2b_1
XFILLER_45_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5460_ _6281_/A _7553_/B vssd1 vssd1 vccd1 vccd1 _5461_/B sky130_fd_sc_hd__nand2_1
X_4411_ _4735_/A vssd1 vssd1 vccd1 vccd1 _4670_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5391_ _5705_/A _5426_/A vssd1 vssd1 vccd1 vccd1 _5562_/A sky130_fd_sc_hd__nor2_1
X_7130_ _7153_/A _7111_/B _7129_/X vssd1 vssd1 vccd1 vccd1 _7139_/A sky130_fd_sc_hd__o21a_1
X_4342_ _4345_/A vssd1 vssd1 vccd1 vccd1 _4342_/Y sky130_fd_sc_hd__inv_2
X_7061_ _7114_/A _7114_/B vssd1 vssd1 vccd1 vccd1 _7064_/B sky130_fd_sc_hd__or2_1
X_4273_ _4277_/A vssd1 vssd1 vccd1 vccd1 _4273_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6012_ _5954_/A _6012_/B vssd1 vssd1 vccd1 vccd1 _6042_/A sky130_fd_sc_hd__and2b_1
.ends

