magic
tech sky130A
magscale 1 2
timestamp 1647759500
<< obsli1 >>
rect 1104 527 58880 53329
<< obsm1 >>
rect 566 280 59418 53848
<< metal2 >>
rect 542 55200 654 56000
rect 1646 55200 1758 56000
rect 2750 55200 2862 56000
rect 3854 55200 3966 56000
rect 4958 55200 5070 56000
rect 6062 55200 6174 56000
rect 7166 55200 7278 56000
rect 8270 55200 8382 56000
rect 9374 55200 9486 56000
rect 10478 55200 10590 56000
rect 11582 55200 11694 56000
rect 12686 55200 12798 56000
rect 13790 55200 13902 56000
rect 14894 55200 15006 56000
rect 16090 55200 16202 56000
rect 17194 55200 17306 56000
rect 18298 55200 18410 56000
rect 19402 55200 19514 56000
rect 20506 55200 20618 56000
rect 21610 55200 21722 56000
rect 22714 55200 22826 56000
rect 23818 55200 23930 56000
rect 24922 55200 25034 56000
rect 26026 55200 26138 56000
rect 27130 55200 27242 56000
rect 28234 55200 28346 56000
rect 29338 55200 29450 56000
rect 30534 55200 30646 56000
rect 31638 55200 31750 56000
rect 32742 55200 32854 56000
rect 33846 55200 33958 56000
rect 34950 55200 35062 56000
rect 36054 55200 36166 56000
rect 37158 55200 37270 56000
rect 38262 55200 38374 56000
rect 39366 55200 39478 56000
rect 40470 55200 40582 56000
rect 41574 55200 41686 56000
rect 42678 55200 42790 56000
rect 43782 55200 43894 56000
rect 44886 55200 44998 56000
rect 46082 55200 46194 56000
rect 47186 55200 47298 56000
rect 48290 55200 48402 56000
rect 49394 55200 49506 56000
rect 50498 55200 50610 56000
rect 51602 55200 51714 56000
rect 52706 55200 52818 56000
rect 53810 55200 53922 56000
rect 54914 55200 55026 56000
rect 56018 55200 56130 56000
rect 57122 55200 57234 56000
rect 58226 55200 58338 56000
rect 59330 55200 59442 56000
rect 3670 0 3782 800
rect 11122 0 11234 800
rect 18666 0 18778 800
rect 26118 0 26230 800
rect 33662 0 33774 800
rect 41114 0 41226 800
rect 48658 0 48770 800
rect 56110 0 56222 800
<< obsm2 >>
rect 710 55144 1590 55593
rect 1814 55144 2694 55593
rect 2918 55144 3798 55593
rect 4022 55144 4902 55593
rect 5126 55144 6006 55593
rect 6230 55144 7110 55593
rect 7334 55144 8214 55593
rect 8438 55144 9318 55593
rect 9542 55144 10422 55593
rect 10646 55144 11526 55593
rect 11750 55144 12630 55593
rect 12854 55144 13734 55593
rect 13958 55144 14838 55593
rect 15062 55144 16034 55593
rect 16258 55144 17138 55593
rect 17362 55144 18242 55593
rect 18466 55144 19346 55593
rect 19570 55144 20450 55593
rect 20674 55144 21554 55593
rect 21778 55144 22658 55593
rect 22882 55144 23762 55593
rect 23986 55144 24866 55593
rect 25090 55144 25970 55593
rect 26194 55144 27074 55593
rect 27298 55144 28178 55593
rect 28402 55144 29282 55593
rect 29506 55144 30478 55593
rect 30702 55144 31582 55593
rect 31806 55144 32686 55593
rect 32910 55144 33790 55593
rect 34014 55144 34894 55593
rect 35118 55144 35998 55593
rect 36222 55144 37102 55593
rect 37326 55144 38206 55593
rect 38430 55144 39310 55593
rect 39534 55144 40414 55593
rect 40638 55144 41518 55593
rect 41742 55144 42622 55593
rect 42846 55144 43726 55593
rect 43950 55144 44830 55593
rect 45054 55144 46026 55593
rect 46250 55144 47130 55593
rect 47354 55144 48234 55593
rect 48458 55144 49338 55593
rect 49562 55144 50442 55593
rect 50666 55144 51546 55593
rect 51770 55144 52650 55593
rect 52874 55144 53754 55593
rect 53978 55144 54858 55593
rect 55082 55144 55962 55593
rect 56186 55144 57066 55593
rect 57290 55144 58170 55593
rect 58394 55144 59274 55593
rect 572 856 59412 55144
rect 572 274 3614 856
rect 3838 274 11066 856
rect 11290 274 18610 856
rect 18834 274 26062 856
rect 26286 274 33606 856
rect 33830 274 41058 856
rect 41282 274 48602 856
rect 48826 274 56054 856
rect 56278 274 59412 856
<< metal3 >>
rect 0 55436 800 55676
rect 59200 55436 60000 55676
rect 0 54620 800 54860
rect 59200 54756 60000 54996
rect 0 53804 800 54044
rect 59200 54076 60000 54316
rect 59200 53396 60000 53636
rect 0 52988 800 53228
rect 59200 52716 60000 52956
rect 0 52172 800 52412
rect 59200 52036 60000 52276
rect 0 51356 800 51596
rect 59200 51356 60000 51596
rect 0 50540 800 50780
rect 59200 50676 60000 50916
rect 0 49724 800 49964
rect 59200 49996 60000 50236
rect 59200 49316 60000 49556
rect 0 48908 800 49148
rect 59200 48636 60000 48876
rect 0 48092 800 48332
rect 59200 47820 60000 48060
rect 0 47276 800 47516
rect 59200 47140 60000 47380
rect 0 46460 800 46700
rect 59200 46460 60000 46700
rect 0 45644 800 45884
rect 59200 45780 60000 46020
rect 0 44828 800 45068
rect 59200 45100 60000 45340
rect 59200 44420 60000 44660
rect 0 44012 800 44252
rect 59200 43740 60000 43980
rect 0 43196 800 43436
rect 59200 43060 60000 43300
rect 0 42380 800 42620
rect 59200 42380 60000 42620
rect 0 41564 800 41804
rect 59200 41700 60000 41940
rect 0 40748 800 40988
rect 59200 41020 60000 41260
rect 59200 40340 60000 40580
rect 0 39932 800 40172
rect 59200 39524 60000 39764
rect 0 39116 800 39356
rect 59200 38844 60000 39084
rect 0 38300 800 38540
rect 59200 38164 60000 38404
rect 0 37484 800 37724
rect 59200 37484 60000 37724
rect 0 36668 800 36908
rect 59200 36804 60000 37044
rect 0 35852 800 36092
rect 59200 36124 60000 36364
rect 59200 35444 60000 35684
rect 0 35036 800 35276
rect 59200 34764 60000 35004
rect 0 34220 800 34460
rect 59200 34084 60000 34324
rect 0 33404 800 33644
rect 59200 33404 60000 33644
rect 0 32588 800 32828
rect 59200 32724 60000 32964
rect 0 31772 800 32012
rect 59200 31908 60000 32148
rect 0 30956 800 31196
rect 59200 31228 60000 31468
rect 59200 30548 60000 30788
rect 0 30140 800 30380
rect 59200 29868 60000 30108
rect 0 29324 800 29564
rect 59200 29188 60000 29428
rect 0 28508 800 28748
rect 59200 28508 60000 28748
rect 0 27828 800 28068
rect 59200 27828 60000 28068
rect 0 27012 800 27252
rect 59200 27148 60000 27388
rect 0 26196 800 26436
rect 59200 26468 60000 26708
rect 59200 25788 60000 26028
rect 0 25380 800 25620
rect 59200 25108 60000 25348
rect 0 24564 800 24804
rect 59200 24428 60000 24668
rect 0 23748 800 23988
rect 59200 23612 60000 23852
rect 0 22932 800 23172
rect 59200 22932 60000 23172
rect 0 22116 800 22356
rect 59200 22252 60000 22492
rect 0 21300 800 21540
rect 59200 21572 60000 21812
rect 59200 20892 60000 21132
rect 0 20484 800 20724
rect 59200 20212 60000 20452
rect 0 19668 800 19908
rect 59200 19532 60000 19772
rect 0 18852 800 19092
rect 59200 18852 60000 19092
rect 0 18036 800 18276
rect 59200 18172 60000 18412
rect 0 17220 800 17460
rect 59200 17492 60000 17732
rect 59200 16812 60000 17052
rect 0 16404 800 16644
rect 59200 15996 60000 16236
rect 0 15588 800 15828
rect 59200 15316 60000 15556
rect 0 14772 800 15012
rect 59200 14636 60000 14876
rect 0 13956 800 14196
rect 59200 13956 60000 14196
rect 0 13140 800 13380
rect 59200 13276 60000 13516
rect 0 12324 800 12564
rect 59200 12596 60000 12836
rect 59200 11916 60000 12156
rect 0 11508 800 11748
rect 59200 11236 60000 11476
rect 0 10692 800 10932
rect 59200 10556 60000 10796
rect 0 9876 800 10116
rect 59200 9876 60000 10116
rect 0 9060 800 9300
rect 59200 9196 60000 9436
rect 0 8244 800 8484
rect 59200 8516 60000 8756
rect 0 7428 800 7668
rect 59200 7700 60000 7940
rect 59200 7020 60000 7260
rect 0 6612 800 6852
rect 59200 6340 60000 6580
rect 0 5796 800 6036
rect 59200 5660 60000 5900
rect 0 4980 800 5220
rect 59200 4980 60000 5220
rect 0 4164 800 4404
rect 59200 4300 60000 4540
rect 0 3348 800 3588
rect 59200 3620 60000 3860
rect 59200 2940 60000 3180
rect 0 2532 800 2772
rect 59200 2260 60000 2500
rect 0 1716 800 1956
rect 59200 1580 60000 1820
rect 0 900 800 1140
rect 59200 900 60000 1140
rect 0 220 800 460
rect 59200 220 60000 460
<< obsm3 >>
rect 880 55356 59120 55589
rect 800 55076 59200 55356
rect 800 54940 59120 55076
rect 880 54676 59120 54940
rect 880 54540 59200 54676
rect 800 54396 59200 54540
rect 800 54124 59120 54396
rect 880 53996 59120 54124
rect 880 53724 59200 53996
rect 800 53716 59200 53724
rect 800 53316 59120 53716
rect 800 53308 59200 53316
rect 880 53036 59200 53308
rect 880 52908 59120 53036
rect 800 52636 59120 52908
rect 800 52492 59200 52636
rect 880 52356 59200 52492
rect 880 52092 59120 52356
rect 800 51956 59120 52092
rect 800 51676 59200 51956
rect 880 51276 59120 51676
rect 800 50996 59200 51276
rect 800 50860 59120 50996
rect 880 50596 59120 50860
rect 880 50460 59200 50596
rect 800 50316 59200 50460
rect 800 50044 59120 50316
rect 880 49916 59120 50044
rect 880 49644 59200 49916
rect 800 49636 59200 49644
rect 800 49236 59120 49636
rect 800 49228 59200 49236
rect 880 48956 59200 49228
rect 880 48828 59120 48956
rect 800 48556 59120 48828
rect 800 48412 59200 48556
rect 880 48140 59200 48412
rect 880 48012 59120 48140
rect 800 47740 59120 48012
rect 800 47596 59200 47740
rect 880 47460 59200 47596
rect 880 47196 59120 47460
rect 800 47060 59120 47196
rect 800 46780 59200 47060
rect 880 46380 59120 46780
rect 800 46100 59200 46380
rect 800 45964 59120 46100
rect 880 45700 59120 45964
rect 880 45564 59200 45700
rect 800 45420 59200 45564
rect 800 45148 59120 45420
rect 880 45020 59120 45148
rect 880 44748 59200 45020
rect 800 44740 59200 44748
rect 800 44340 59120 44740
rect 800 44332 59200 44340
rect 880 44060 59200 44332
rect 880 43932 59120 44060
rect 800 43660 59120 43932
rect 800 43516 59200 43660
rect 880 43380 59200 43516
rect 880 43116 59120 43380
rect 800 42980 59120 43116
rect 800 42700 59200 42980
rect 880 42300 59120 42700
rect 800 42020 59200 42300
rect 800 41884 59120 42020
rect 880 41620 59120 41884
rect 880 41484 59200 41620
rect 800 41340 59200 41484
rect 800 41068 59120 41340
rect 880 40940 59120 41068
rect 880 40668 59200 40940
rect 800 40660 59200 40668
rect 800 40260 59120 40660
rect 800 40252 59200 40260
rect 880 39852 59200 40252
rect 800 39844 59200 39852
rect 800 39444 59120 39844
rect 800 39436 59200 39444
rect 880 39164 59200 39436
rect 880 39036 59120 39164
rect 800 38764 59120 39036
rect 800 38620 59200 38764
rect 880 38484 59200 38620
rect 880 38220 59120 38484
rect 800 38084 59120 38220
rect 800 37804 59200 38084
rect 880 37404 59120 37804
rect 800 37124 59200 37404
rect 800 36988 59120 37124
rect 880 36724 59120 36988
rect 880 36588 59200 36724
rect 800 36444 59200 36588
rect 800 36172 59120 36444
rect 880 36044 59120 36172
rect 880 35772 59200 36044
rect 800 35764 59200 35772
rect 800 35364 59120 35764
rect 800 35356 59200 35364
rect 880 35084 59200 35356
rect 880 34956 59120 35084
rect 800 34684 59120 34956
rect 800 34540 59200 34684
rect 880 34404 59200 34540
rect 880 34140 59120 34404
rect 800 34004 59120 34140
rect 800 33724 59200 34004
rect 880 33324 59120 33724
rect 800 33044 59200 33324
rect 800 32908 59120 33044
rect 880 32644 59120 32908
rect 880 32508 59200 32644
rect 800 32228 59200 32508
rect 800 32092 59120 32228
rect 880 31828 59120 32092
rect 880 31692 59200 31828
rect 800 31548 59200 31692
rect 800 31276 59120 31548
rect 880 31148 59120 31276
rect 880 30876 59200 31148
rect 800 30868 59200 30876
rect 800 30468 59120 30868
rect 800 30460 59200 30468
rect 880 30188 59200 30460
rect 880 30060 59120 30188
rect 800 29788 59120 30060
rect 800 29644 59200 29788
rect 880 29508 59200 29644
rect 880 29244 59120 29508
rect 800 29108 59120 29244
rect 800 28828 59200 29108
rect 880 28428 59120 28828
rect 800 28148 59200 28428
rect 880 27748 59120 28148
rect 800 27468 59200 27748
rect 800 27332 59120 27468
rect 880 27068 59120 27332
rect 880 26932 59200 27068
rect 800 26788 59200 26932
rect 800 26516 59120 26788
rect 880 26388 59120 26516
rect 880 26116 59200 26388
rect 800 26108 59200 26116
rect 800 25708 59120 26108
rect 800 25700 59200 25708
rect 880 25428 59200 25700
rect 880 25300 59120 25428
rect 800 25028 59120 25300
rect 800 24884 59200 25028
rect 880 24748 59200 24884
rect 880 24484 59120 24748
rect 800 24348 59120 24484
rect 800 24068 59200 24348
rect 880 23932 59200 24068
rect 880 23668 59120 23932
rect 800 23532 59120 23668
rect 800 23252 59200 23532
rect 880 22852 59120 23252
rect 800 22572 59200 22852
rect 800 22436 59120 22572
rect 880 22172 59120 22436
rect 880 22036 59200 22172
rect 800 21892 59200 22036
rect 800 21620 59120 21892
rect 880 21492 59120 21620
rect 880 21220 59200 21492
rect 800 21212 59200 21220
rect 800 20812 59120 21212
rect 800 20804 59200 20812
rect 880 20532 59200 20804
rect 880 20404 59120 20532
rect 800 20132 59120 20404
rect 800 19988 59200 20132
rect 880 19852 59200 19988
rect 880 19588 59120 19852
rect 800 19452 59120 19588
rect 800 19172 59200 19452
rect 880 18772 59120 19172
rect 800 18492 59200 18772
rect 800 18356 59120 18492
rect 880 18092 59120 18356
rect 880 17956 59200 18092
rect 800 17812 59200 17956
rect 800 17540 59120 17812
rect 880 17412 59120 17540
rect 880 17140 59200 17412
rect 800 17132 59200 17140
rect 800 16732 59120 17132
rect 800 16724 59200 16732
rect 880 16324 59200 16724
rect 800 16316 59200 16324
rect 800 15916 59120 16316
rect 800 15908 59200 15916
rect 880 15636 59200 15908
rect 880 15508 59120 15636
rect 800 15236 59120 15508
rect 800 15092 59200 15236
rect 880 14956 59200 15092
rect 880 14692 59120 14956
rect 800 14556 59120 14692
rect 800 14276 59200 14556
rect 880 13876 59120 14276
rect 800 13596 59200 13876
rect 800 13460 59120 13596
rect 880 13196 59120 13460
rect 880 13060 59200 13196
rect 800 12916 59200 13060
rect 800 12644 59120 12916
rect 880 12516 59120 12644
rect 880 12244 59200 12516
rect 800 12236 59200 12244
rect 800 11836 59120 12236
rect 800 11828 59200 11836
rect 880 11556 59200 11828
rect 880 11428 59120 11556
rect 800 11156 59120 11428
rect 800 11012 59200 11156
rect 880 10876 59200 11012
rect 880 10612 59120 10876
rect 800 10476 59120 10612
rect 800 10196 59200 10476
rect 880 9796 59120 10196
rect 800 9516 59200 9796
rect 800 9380 59120 9516
rect 880 9116 59120 9380
rect 880 8980 59200 9116
rect 800 8836 59200 8980
rect 800 8564 59120 8836
rect 880 8436 59120 8564
rect 880 8164 59200 8436
rect 800 8020 59200 8164
rect 800 7748 59120 8020
rect 880 7620 59120 7748
rect 880 7348 59200 7620
rect 800 7340 59200 7348
rect 800 6940 59120 7340
rect 800 6932 59200 6940
rect 880 6660 59200 6932
rect 880 6532 59120 6660
rect 800 6260 59120 6532
rect 800 6116 59200 6260
rect 880 5980 59200 6116
rect 880 5716 59120 5980
rect 800 5580 59120 5716
rect 800 5300 59200 5580
rect 880 4900 59120 5300
rect 800 4620 59200 4900
rect 800 4484 59120 4620
rect 880 4220 59120 4484
rect 880 4084 59200 4220
rect 800 3940 59200 4084
rect 800 3668 59120 3940
rect 880 3540 59120 3668
rect 880 3268 59200 3540
rect 800 3260 59200 3268
rect 800 2860 59120 3260
rect 800 2852 59200 2860
rect 880 2580 59200 2852
rect 880 2452 59120 2580
rect 800 2180 59120 2452
rect 800 2036 59200 2180
rect 880 1900 59200 2036
rect 880 1636 59120 1900
rect 800 1500 59120 1636
rect 800 1220 59200 1500
rect 880 820 59120 1220
rect 800 540 59200 820
rect 880 511 59120 540
<< metal4 >>
rect 4208 496 4528 53360
rect 19568 496 19888 53360
rect 34928 496 35248 53360
rect 50288 496 50608 53360
<< obsm4 >>
rect 6867 579 19488 46477
rect 19968 579 34848 46477
rect 35328 579 39133 46477
<< labels >>
rlabel metal2 s 542 55200 654 56000 6 active
port 1 nsew signal input
rlabel metal2 s 2750 55200 2862 56000 6 io_in[0]
port 2 nsew signal input
rlabel metal2 s 13790 55200 13902 56000 6 io_in[10]
port 3 nsew signal input
rlabel metal2 s 14894 55200 15006 56000 6 io_in[11]
port 4 nsew signal input
rlabel metal2 s 16090 55200 16202 56000 6 io_in[12]
port 5 nsew signal input
rlabel metal2 s 17194 55200 17306 56000 6 io_in[13]
port 6 nsew signal input
rlabel metal2 s 18298 55200 18410 56000 6 io_in[14]
port 7 nsew signal input
rlabel metal2 s 19402 55200 19514 56000 6 io_in[15]
port 8 nsew signal input
rlabel metal2 s 20506 55200 20618 56000 6 io_in[16]
port 9 nsew signal input
rlabel metal2 s 21610 55200 21722 56000 6 io_in[17]
port 10 nsew signal input
rlabel metal2 s 22714 55200 22826 56000 6 io_in[18]
port 11 nsew signal input
rlabel metal2 s 23818 55200 23930 56000 6 io_in[19]
port 12 nsew signal input
rlabel metal2 s 3854 55200 3966 56000 6 io_in[1]
port 13 nsew signal input
rlabel metal2 s 24922 55200 25034 56000 6 io_in[20]
port 14 nsew signal input
rlabel metal2 s 26026 55200 26138 56000 6 io_in[21]
port 15 nsew signal input
rlabel metal2 s 27130 55200 27242 56000 6 io_in[22]
port 16 nsew signal input
rlabel metal2 s 28234 55200 28346 56000 6 io_in[23]
port 17 nsew signal input
rlabel metal2 s 29338 55200 29450 56000 6 io_in[24]
port 18 nsew signal input
rlabel metal2 s 30534 55200 30646 56000 6 io_in[25]
port 19 nsew signal input
rlabel metal2 s 31638 55200 31750 56000 6 io_in[26]
port 20 nsew signal input
rlabel metal2 s 32742 55200 32854 56000 6 io_in[27]
port 21 nsew signal input
rlabel metal2 s 33846 55200 33958 56000 6 io_in[28]
port 22 nsew signal input
rlabel metal2 s 34950 55200 35062 56000 6 io_in[29]
port 23 nsew signal input
rlabel metal2 s 4958 55200 5070 56000 6 io_in[2]
port 24 nsew signal input
rlabel metal2 s 36054 55200 36166 56000 6 io_in[30]
port 25 nsew signal input
rlabel metal2 s 37158 55200 37270 56000 6 io_in[31]
port 26 nsew signal input
rlabel metal2 s 38262 55200 38374 56000 6 io_in[32]
port 27 nsew signal input
rlabel metal2 s 39366 55200 39478 56000 6 io_in[33]
port 28 nsew signal input
rlabel metal2 s 40470 55200 40582 56000 6 io_in[34]
port 29 nsew signal input
rlabel metal2 s 41574 55200 41686 56000 6 io_in[35]
port 30 nsew signal input
rlabel metal2 s 42678 55200 42790 56000 6 io_in[36]
port 31 nsew signal input
rlabel metal2 s 43782 55200 43894 56000 6 io_in[37]
port 32 nsew signal input
rlabel metal2 s 6062 55200 6174 56000 6 io_in[3]
port 33 nsew signal input
rlabel metal2 s 7166 55200 7278 56000 6 io_in[4]
port 34 nsew signal input
rlabel metal2 s 8270 55200 8382 56000 6 io_in[5]
port 35 nsew signal input
rlabel metal2 s 9374 55200 9486 56000 6 io_in[6]
port 36 nsew signal input
rlabel metal2 s 10478 55200 10590 56000 6 io_in[7]
port 37 nsew signal input
rlabel metal2 s 11582 55200 11694 56000 6 io_in[8]
port 38 nsew signal input
rlabel metal2 s 12686 55200 12798 56000 6 io_in[9]
port 39 nsew signal input
rlabel metal3 s 59200 22252 60000 22492 6 io_oeb[0]
port 40 nsew signal output
rlabel metal3 s 59200 29188 60000 29428 6 io_oeb[10]
port 41 nsew signal output
rlabel metal3 s 59200 29868 60000 30108 6 io_oeb[11]
port 42 nsew signal output
rlabel metal3 s 59200 30548 60000 30788 6 io_oeb[12]
port 43 nsew signal output
rlabel metal3 s 59200 31228 60000 31468 6 io_oeb[13]
port 44 nsew signal output
rlabel metal3 s 59200 31908 60000 32148 6 io_oeb[14]
port 45 nsew signal output
rlabel metal3 s 59200 32724 60000 32964 6 io_oeb[15]
port 46 nsew signal output
rlabel metal3 s 59200 33404 60000 33644 6 io_oeb[16]
port 47 nsew signal output
rlabel metal3 s 59200 34084 60000 34324 6 io_oeb[17]
port 48 nsew signal output
rlabel metal3 s 59200 34764 60000 35004 6 io_oeb[18]
port 49 nsew signal output
rlabel metal3 s 59200 35444 60000 35684 6 io_oeb[19]
port 50 nsew signal output
rlabel metal3 s 59200 22932 60000 23172 6 io_oeb[1]
port 51 nsew signal output
rlabel metal3 s 59200 36124 60000 36364 6 io_oeb[20]
port 52 nsew signal output
rlabel metal3 s 59200 36804 60000 37044 6 io_oeb[21]
port 53 nsew signal output
rlabel metal3 s 59200 37484 60000 37724 6 io_oeb[22]
port 54 nsew signal output
rlabel metal3 s 59200 38164 60000 38404 6 io_oeb[23]
port 55 nsew signal output
rlabel metal3 s 59200 38844 60000 39084 6 io_oeb[24]
port 56 nsew signal output
rlabel metal3 s 59200 39524 60000 39764 6 io_oeb[25]
port 57 nsew signal output
rlabel metal3 s 59200 40340 60000 40580 6 io_oeb[26]
port 58 nsew signal output
rlabel metal3 s 59200 41020 60000 41260 6 io_oeb[27]
port 59 nsew signal output
rlabel metal3 s 59200 41700 60000 41940 6 io_oeb[28]
port 60 nsew signal output
rlabel metal3 s 59200 42380 60000 42620 6 io_oeb[29]
port 61 nsew signal output
rlabel metal3 s 59200 23612 60000 23852 6 io_oeb[2]
port 62 nsew signal output
rlabel metal3 s 59200 43060 60000 43300 6 io_oeb[30]
port 63 nsew signal output
rlabel metal3 s 59200 43740 60000 43980 6 io_oeb[31]
port 64 nsew signal output
rlabel metal3 s 59200 44420 60000 44660 6 io_oeb[32]
port 65 nsew signal output
rlabel metal3 s 59200 45100 60000 45340 6 io_oeb[33]
port 66 nsew signal output
rlabel metal3 s 59200 45780 60000 46020 6 io_oeb[34]
port 67 nsew signal output
rlabel metal3 s 59200 46460 60000 46700 6 io_oeb[35]
port 68 nsew signal output
rlabel metal3 s 59200 47140 60000 47380 6 io_oeb[36]
port 69 nsew signal output
rlabel metal3 s 59200 47820 60000 48060 6 io_oeb[37]
port 70 nsew signal output
rlabel metal3 s 59200 24428 60000 24668 6 io_oeb[3]
port 71 nsew signal output
rlabel metal3 s 59200 25108 60000 25348 6 io_oeb[4]
port 72 nsew signal output
rlabel metal3 s 59200 25788 60000 26028 6 io_oeb[5]
port 73 nsew signal output
rlabel metal3 s 59200 26468 60000 26708 6 io_oeb[6]
port 74 nsew signal output
rlabel metal3 s 59200 27148 60000 27388 6 io_oeb[7]
port 75 nsew signal output
rlabel metal3 s 59200 27828 60000 28068 6 io_oeb[8]
port 76 nsew signal output
rlabel metal3 s 59200 28508 60000 28748 6 io_oeb[9]
port 77 nsew signal output
rlabel metal3 s 59200 48636 60000 48876 6 io_out[0]
port 78 nsew signal output
rlabel metal3 s 59200 50676 60000 50916 6 io_out[10]
port 79 nsew signal output
rlabel metal3 s 59200 51356 60000 51596 6 io_out[11]
port 80 nsew signal output
rlabel metal2 s 11122 0 11234 800 6 io_out[12]
port 81 nsew signal output
rlabel metal2 s 50498 55200 50610 56000 6 io_out[13]
port 82 nsew signal output
rlabel metal2 s 18666 0 18778 800 6 io_out[14]
port 83 nsew signal output
rlabel metal2 s 26118 0 26230 800 6 io_out[15]
port 84 nsew signal output
rlabel metal2 s 33662 0 33774 800 6 io_out[16]
port 85 nsew signal output
rlabel metal2 s 51602 55200 51714 56000 6 io_out[17]
port 86 nsew signal output
rlabel metal3 s 59200 52036 60000 52276 6 io_out[18]
port 87 nsew signal output
rlabel metal3 s 59200 52716 60000 52956 6 io_out[19]
port 88 nsew signal output
rlabel metal3 s 0 52172 800 52412 6 io_out[1]
port 89 nsew signal output
rlabel metal2 s 52706 55200 52818 56000 6 io_out[20]
port 90 nsew signal output
rlabel metal3 s 0 52988 800 53228 6 io_out[21]
port 91 nsew signal output
rlabel metal3 s 59200 53396 60000 53636 6 io_out[22]
port 92 nsew signal output
rlabel metal2 s 53810 55200 53922 56000 6 io_out[23]
port 93 nsew signal output
rlabel metal3 s 59200 54076 60000 54316 6 io_out[24]
port 94 nsew signal output
rlabel metal3 s 59200 54756 60000 54996 6 io_out[25]
port 95 nsew signal output
rlabel metal3 s 0 53804 800 54044 6 io_out[26]
port 96 nsew signal output
rlabel metal2 s 54914 55200 55026 56000 6 io_out[27]
port 97 nsew signal output
rlabel metal2 s 56018 55200 56130 56000 6 io_out[28]
port 98 nsew signal output
rlabel metal2 s 57122 55200 57234 56000 6 io_out[29]
port 99 nsew signal output
rlabel metal2 s 44886 55200 44998 56000 6 io_out[2]
port 100 nsew signal output
rlabel metal2 s 58226 55200 58338 56000 6 io_out[30]
port 101 nsew signal output
rlabel metal2 s 41114 0 41226 800 6 io_out[31]
port 102 nsew signal output
rlabel metal3 s 59200 55436 60000 55676 6 io_out[32]
port 103 nsew signal output
rlabel metal2 s 48658 0 48770 800 6 io_out[33]
port 104 nsew signal output
rlabel metal2 s 56110 0 56222 800 6 io_out[34]
port 105 nsew signal output
rlabel metal3 s 0 54620 800 54860 6 io_out[35]
port 106 nsew signal output
rlabel metal2 s 59330 55200 59442 56000 6 io_out[36]
port 107 nsew signal output
rlabel metal3 s 0 55436 800 55676 6 io_out[37]
port 108 nsew signal output
rlabel metal2 s 46082 55200 46194 56000 6 io_out[3]
port 109 nsew signal output
rlabel metal2 s 47186 55200 47298 56000 6 io_out[4]
port 110 nsew signal output
rlabel metal2 s 3670 0 3782 800 6 io_out[5]
port 111 nsew signal output
rlabel metal2 s 48290 55200 48402 56000 6 io_out[6]
port 112 nsew signal output
rlabel metal3 s 59200 49316 60000 49556 6 io_out[7]
port 113 nsew signal output
rlabel metal3 s 59200 49996 60000 50236 6 io_out[8]
port 114 nsew signal output
rlabel metal2 s 49394 55200 49506 56000 6 io_out[9]
port 115 nsew signal output
rlabel metal3 s 0 220 800 460 6 la1_data_in[0]
port 116 nsew signal input
rlabel metal3 s 0 8244 800 8484 6 la1_data_in[10]
port 117 nsew signal input
rlabel metal3 s 0 9060 800 9300 6 la1_data_in[11]
port 118 nsew signal input
rlabel metal3 s 0 9876 800 10116 6 la1_data_in[12]
port 119 nsew signal input
rlabel metal3 s 0 10692 800 10932 6 la1_data_in[13]
port 120 nsew signal input
rlabel metal3 s 0 11508 800 11748 6 la1_data_in[14]
port 121 nsew signal input
rlabel metal3 s 0 12324 800 12564 6 la1_data_in[15]
port 122 nsew signal input
rlabel metal3 s 0 13140 800 13380 6 la1_data_in[16]
port 123 nsew signal input
rlabel metal3 s 0 13956 800 14196 6 la1_data_in[17]
port 124 nsew signal input
rlabel metal3 s 0 14772 800 15012 6 la1_data_in[18]
port 125 nsew signal input
rlabel metal3 s 0 15588 800 15828 6 la1_data_in[19]
port 126 nsew signal input
rlabel metal3 s 0 900 800 1140 6 la1_data_in[1]
port 127 nsew signal input
rlabel metal3 s 0 16404 800 16644 6 la1_data_in[20]
port 128 nsew signal input
rlabel metal3 s 0 17220 800 17460 6 la1_data_in[21]
port 129 nsew signal input
rlabel metal3 s 0 18036 800 18276 6 la1_data_in[22]
port 130 nsew signal input
rlabel metal3 s 0 18852 800 19092 6 la1_data_in[23]
port 131 nsew signal input
rlabel metal3 s 0 19668 800 19908 6 la1_data_in[24]
port 132 nsew signal input
rlabel metal3 s 0 20484 800 20724 6 la1_data_in[25]
port 133 nsew signal input
rlabel metal3 s 0 21300 800 21540 6 la1_data_in[26]
port 134 nsew signal input
rlabel metal3 s 0 22116 800 22356 6 la1_data_in[27]
port 135 nsew signal input
rlabel metal3 s 0 22932 800 23172 6 la1_data_in[28]
port 136 nsew signal input
rlabel metal3 s 0 23748 800 23988 6 la1_data_in[29]
port 137 nsew signal input
rlabel metal3 s 0 1716 800 1956 6 la1_data_in[2]
port 138 nsew signal input
rlabel metal3 s 0 24564 800 24804 6 la1_data_in[30]
port 139 nsew signal input
rlabel metal3 s 0 25380 800 25620 6 la1_data_in[31]
port 140 nsew signal input
rlabel metal3 s 0 2532 800 2772 6 la1_data_in[3]
port 141 nsew signal input
rlabel metal3 s 0 3348 800 3588 6 la1_data_in[4]
port 142 nsew signal input
rlabel metal3 s 0 4164 800 4404 6 la1_data_in[5]
port 143 nsew signal input
rlabel metal3 s 0 4980 800 5220 6 la1_data_in[6]
port 144 nsew signal input
rlabel metal3 s 0 5796 800 6036 6 la1_data_in[7]
port 145 nsew signal input
rlabel metal3 s 0 6612 800 6852 6 la1_data_in[8]
port 146 nsew signal input
rlabel metal3 s 0 7428 800 7668 6 la1_data_in[9]
port 147 nsew signal input
rlabel metal3 s 0 26196 800 26436 6 la1_data_out[0]
port 148 nsew signal output
rlabel metal3 s 0 34220 800 34460 6 la1_data_out[10]
port 149 nsew signal output
rlabel metal3 s 0 35036 800 35276 6 la1_data_out[11]
port 150 nsew signal output
rlabel metal3 s 0 35852 800 36092 6 la1_data_out[12]
port 151 nsew signal output
rlabel metal3 s 0 36668 800 36908 6 la1_data_out[13]
port 152 nsew signal output
rlabel metal3 s 0 37484 800 37724 6 la1_data_out[14]
port 153 nsew signal output
rlabel metal3 s 0 38300 800 38540 6 la1_data_out[15]
port 154 nsew signal output
rlabel metal3 s 0 39116 800 39356 6 la1_data_out[16]
port 155 nsew signal output
rlabel metal3 s 0 39932 800 40172 6 la1_data_out[17]
port 156 nsew signal output
rlabel metal3 s 0 40748 800 40988 6 la1_data_out[18]
port 157 nsew signal output
rlabel metal3 s 0 41564 800 41804 6 la1_data_out[19]
port 158 nsew signal output
rlabel metal3 s 0 27012 800 27252 6 la1_data_out[1]
port 159 nsew signal output
rlabel metal3 s 0 42380 800 42620 6 la1_data_out[20]
port 160 nsew signal output
rlabel metal3 s 0 43196 800 43436 6 la1_data_out[21]
port 161 nsew signal output
rlabel metal3 s 0 44012 800 44252 6 la1_data_out[22]
port 162 nsew signal output
rlabel metal3 s 0 44828 800 45068 6 la1_data_out[23]
port 163 nsew signal output
rlabel metal3 s 0 45644 800 45884 6 la1_data_out[24]
port 164 nsew signal output
rlabel metal3 s 0 46460 800 46700 6 la1_data_out[25]
port 165 nsew signal output
rlabel metal3 s 0 47276 800 47516 6 la1_data_out[26]
port 166 nsew signal output
rlabel metal3 s 0 48092 800 48332 6 la1_data_out[27]
port 167 nsew signal output
rlabel metal3 s 0 48908 800 49148 6 la1_data_out[28]
port 168 nsew signal output
rlabel metal3 s 0 49724 800 49964 6 la1_data_out[29]
port 169 nsew signal output
rlabel metal3 s 0 27828 800 28068 6 la1_data_out[2]
port 170 nsew signal output
rlabel metal3 s 0 50540 800 50780 6 la1_data_out[30]
port 171 nsew signal output
rlabel metal3 s 0 51356 800 51596 6 la1_data_out[31]
port 172 nsew signal output
rlabel metal3 s 0 28508 800 28748 6 la1_data_out[3]
port 173 nsew signal output
rlabel metal3 s 0 29324 800 29564 6 la1_data_out[4]
port 174 nsew signal output
rlabel metal3 s 0 30140 800 30380 6 la1_data_out[5]
port 175 nsew signal output
rlabel metal3 s 0 30956 800 31196 6 la1_data_out[6]
port 176 nsew signal output
rlabel metal3 s 0 31772 800 32012 6 la1_data_out[7]
port 177 nsew signal output
rlabel metal3 s 0 32588 800 32828 6 la1_data_out[8]
port 178 nsew signal output
rlabel metal3 s 0 33404 800 33644 6 la1_data_out[9]
port 179 nsew signal output
rlabel metal3 s 59200 220 60000 460 6 la1_oenb[0]
port 180 nsew signal input
rlabel metal3 s 59200 7020 60000 7260 6 la1_oenb[10]
port 181 nsew signal input
rlabel metal3 s 59200 7700 60000 7940 6 la1_oenb[11]
port 182 nsew signal input
rlabel metal3 s 59200 8516 60000 8756 6 la1_oenb[12]
port 183 nsew signal input
rlabel metal3 s 59200 9196 60000 9436 6 la1_oenb[13]
port 184 nsew signal input
rlabel metal3 s 59200 9876 60000 10116 6 la1_oenb[14]
port 185 nsew signal input
rlabel metal3 s 59200 10556 60000 10796 6 la1_oenb[15]
port 186 nsew signal input
rlabel metal3 s 59200 11236 60000 11476 6 la1_oenb[16]
port 187 nsew signal input
rlabel metal3 s 59200 11916 60000 12156 6 la1_oenb[17]
port 188 nsew signal input
rlabel metal3 s 59200 12596 60000 12836 6 la1_oenb[18]
port 189 nsew signal input
rlabel metal3 s 59200 13276 60000 13516 6 la1_oenb[19]
port 190 nsew signal input
rlabel metal3 s 59200 900 60000 1140 6 la1_oenb[1]
port 191 nsew signal input
rlabel metal3 s 59200 13956 60000 14196 6 la1_oenb[20]
port 192 nsew signal input
rlabel metal3 s 59200 14636 60000 14876 6 la1_oenb[21]
port 193 nsew signal input
rlabel metal3 s 59200 15316 60000 15556 6 la1_oenb[22]
port 194 nsew signal input
rlabel metal3 s 59200 15996 60000 16236 6 la1_oenb[23]
port 195 nsew signal input
rlabel metal3 s 59200 16812 60000 17052 6 la1_oenb[24]
port 196 nsew signal input
rlabel metal3 s 59200 17492 60000 17732 6 la1_oenb[25]
port 197 nsew signal input
rlabel metal3 s 59200 18172 60000 18412 6 la1_oenb[26]
port 198 nsew signal input
rlabel metal3 s 59200 18852 60000 19092 6 la1_oenb[27]
port 199 nsew signal input
rlabel metal3 s 59200 19532 60000 19772 6 la1_oenb[28]
port 200 nsew signal input
rlabel metal3 s 59200 20212 60000 20452 6 la1_oenb[29]
port 201 nsew signal input
rlabel metal3 s 59200 1580 60000 1820 6 la1_oenb[2]
port 202 nsew signal input
rlabel metal3 s 59200 20892 60000 21132 6 la1_oenb[30]
port 203 nsew signal input
rlabel metal3 s 59200 21572 60000 21812 6 la1_oenb[31]
port 204 nsew signal input
rlabel metal3 s 59200 2260 60000 2500 6 la1_oenb[3]
port 205 nsew signal input
rlabel metal3 s 59200 2940 60000 3180 6 la1_oenb[4]
port 206 nsew signal input
rlabel metal3 s 59200 3620 60000 3860 6 la1_oenb[5]
port 207 nsew signal input
rlabel metal3 s 59200 4300 60000 4540 6 la1_oenb[6]
port 208 nsew signal input
rlabel metal3 s 59200 4980 60000 5220 6 la1_oenb[7]
port 209 nsew signal input
rlabel metal3 s 59200 5660 60000 5900 6 la1_oenb[8]
port 210 nsew signal input
rlabel metal3 s 59200 6340 60000 6580 6 la1_oenb[9]
port 211 nsew signal input
rlabel metal4 s 4208 496 4528 53360 6 vccd1
port 212 nsew power input
rlabel metal4 s 34928 496 35248 53360 6 vccd1
port 212 nsew power input
rlabel metal4 s 19568 496 19888 53360 6 vssd1
port 213 nsew ground input
rlabel metal4 s 50288 496 50608 53360 6 vssd1
port 213 nsew ground input
rlabel metal2 s 1646 55200 1758 56000 6 wb_clk_i
port 214 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 60000 56000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 12595880
string GDS_FILE /openlane/designs/wrapped-vgademo-on-fpga/runs/RUN_2022.03.20_06.53.13/results/finishing/wrapped_vgademo_on_fpga.magic.gds
string GDS_START 1116876
<< end >>

